module RegsRouter( // @[:@3.2]
  input  [2:0]  io_selector, // @[:@6.4]
  input  [31:0] io_input_regs_0_ra, // @[:@6.4]
  input  [31:0] io_input_regs_0_sp, // @[:@6.4]
  input  [31:0] io_input_regs_0_gp, // @[:@6.4]
  input  [31:0] io_input_regs_0_tp, // @[:@6.4]
  input  [31:0] io_input_regs_0_t0, // @[:@6.4]
  input  [31:0] io_input_regs_0_t1, // @[:@6.4]
  input  [31:0] io_input_regs_0_t2, // @[:@6.4]
  input  [31:0] io_input_regs_0_fp, // @[:@6.4]
  input  [31:0] io_input_regs_0_s1, // @[:@6.4]
  input  [31:0] io_input_regs_0_a0, // @[:@6.4]
  input  [31:0] io_input_regs_0_a1, // @[:@6.4]
  input  [31:0] io_input_regs_0_a2, // @[:@6.4]
  input  [31:0] io_input_regs_0_a3, // @[:@6.4]
  input  [31:0] io_input_regs_0_a4, // @[:@6.4]
  input  [31:0] io_input_regs_0_a5, // @[:@6.4]
  input  [31:0] io_input_regs_0_a6, // @[:@6.4]
  input  [31:0] io_input_regs_0_a7, // @[:@6.4]
  input  [31:0] io_input_regs_0_s2, // @[:@6.4]
  input  [31:0] io_input_regs_0_s3, // @[:@6.4]
  input  [31:0] io_input_regs_0_s4, // @[:@6.4]
  input  [31:0] io_input_regs_0_s5, // @[:@6.4]
  input  [31:0] io_input_regs_0_s6, // @[:@6.4]
  input  [31:0] io_input_regs_0_s7, // @[:@6.4]
  input  [31:0] io_input_regs_0_s8, // @[:@6.4]
  input  [31:0] io_input_regs_0_s9, // @[:@6.4]
  input  [31:0] io_input_regs_0_s10, // @[:@6.4]
  input  [31:0] io_input_regs_0_s11, // @[:@6.4]
  input  [31:0] io_input_regs_0_t3, // @[:@6.4]
  input  [31:0] io_input_regs_0_t4, // @[:@6.4]
  input  [31:0] io_input_regs_0_t5, // @[:@6.4]
  input  [31:0] io_input_regs_0_t6, // @[:@6.4]
  input  [31:0] io_input_regs_0_pc, // @[:@6.4]
  input         io_input_regs_0_interrupt, // @[:@6.4]
  input  [31:0] io_input_regs_0_interrupt_cause, // @[:@6.4]
  input  [31:0] io_input_regs_0_time, // @[:@6.4]
  input         io_input_regs_0_debug, // @[:@6.4]
  input  [31:0] io_input_regs_0_isa, // @[:@6.4]
  input         io_input_regs_0_sd, // @[:@6.4]
  input         io_input_regs_0_sd_rv32, // @[:@6.4]
  input  [31:0] io_input_regs_0_mpp, // @[:@6.4]
  input         io_input_regs_0_spp, // @[:@6.4]
  input         io_input_regs_0_mpie, // @[:@6.4]
  input         io_input_regs_0_mie, // @[:@6.4]
  input  [31:0] io_input_regs_0_evec, // @[:@6.4]
  input  [31:0] io_input_regs_1_ra, // @[:@6.4]
  input  [31:0] io_input_regs_1_sp, // @[:@6.4]
  input  [31:0] io_input_regs_1_gp, // @[:@6.4]
  input  [31:0] io_input_regs_1_tp, // @[:@6.4]
  input  [31:0] io_input_regs_1_t0, // @[:@6.4]
  input  [31:0] io_input_regs_1_t1, // @[:@6.4]
  input  [31:0] io_input_regs_1_t2, // @[:@6.4]
  input  [31:0] io_input_regs_1_fp, // @[:@6.4]
  input  [31:0] io_input_regs_1_s1, // @[:@6.4]
  input  [31:0] io_input_regs_1_a0, // @[:@6.4]
  input  [31:0] io_input_regs_1_a1, // @[:@6.4]
  input  [31:0] io_input_regs_1_a2, // @[:@6.4]
  input  [31:0] io_input_regs_1_a3, // @[:@6.4]
  input  [31:0] io_input_regs_1_a4, // @[:@6.4]
  input  [31:0] io_input_regs_1_a5, // @[:@6.4]
  input  [31:0] io_input_regs_1_a6, // @[:@6.4]
  input  [31:0] io_input_regs_1_a7, // @[:@6.4]
  input  [31:0] io_input_regs_1_s2, // @[:@6.4]
  input  [31:0] io_input_regs_1_s3, // @[:@6.4]
  input  [31:0] io_input_regs_1_s4, // @[:@6.4]
  input  [31:0] io_input_regs_1_s5, // @[:@6.4]
  input  [31:0] io_input_regs_1_s6, // @[:@6.4]
  input  [31:0] io_input_regs_1_s7, // @[:@6.4]
  input  [31:0] io_input_regs_1_s8, // @[:@6.4]
  input  [31:0] io_input_regs_1_s9, // @[:@6.4]
  input  [31:0] io_input_regs_1_s10, // @[:@6.4]
  input  [31:0] io_input_regs_1_s11, // @[:@6.4]
  input  [31:0] io_input_regs_1_t3, // @[:@6.4]
  input  [31:0] io_input_regs_1_t4, // @[:@6.4]
  input  [31:0] io_input_regs_1_t5, // @[:@6.4]
  input  [31:0] io_input_regs_1_t6, // @[:@6.4]
  input  [31:0] io_input_regs_1_pc, // @[:@6.4]
  input         io_input_regs_1_interrupt, // @[:@6.4]
  input  [31:0] io_input_regs_1_interrupt_cause, // @[:@6.4]
  input  [31:0] io_input_regs_1_time, // @[:@6.4]
  input         io_input_regs_1_debug, // @[:@6.4]
  input  [31:0] io_input_regs_1_isa, // @[:@6.4]
  input         io_input_regs_1_sd, // @[:@6.4]
  input         io_input_regs_1_sd_rv32, // @[:@6.4]
  input  [31:0] io_input_regs_1_mpp, // @[:@6.4]
  input         io_input_regs_1_spp, // @[:@6.4]
  input         io_input_regs_1_mpie, // @[:@6.4]
  input         io_input_regs_1_mie, // @[:@6.4]
  input  [31:0] io_input_regs_1_evec, // @[:@6.4]
  input  [31:0] io_input_regs_2_ra, // @[:@6.4]
  input  [31:0] io_input_regs_2_sp, // @[:@6.4]
  input  [31:0] io_input_regs_2_gp, // @[:@6.4]
  input  [31:0] io_input_regs_2_tp, // @[:@6.4]
  input  [31:0] io_input_regs_2_t0, // @[:@6.4]
  input  [31:0] io_input_regs_2_t1, // @[:@6.4]
  input  [31:0] io_input_regs_2_t2, // @[:@6.4]
  input  [31:0] io_input_regs_2_fp, // @[:@6.4]
  input  [31:0] io_input_regs_2_s1, // @[:@6.4]
  input  [31:0] io_input_regs_2_a0, // @[:@6.4]
  input  [31:0] io_input_regs_2_a1, // @[:@6.4]
  input  [31:0] io_input_regs_2_a2, // @[:@6.4]
  input  [31:0] io_input_regs_2_a3, // @[:@6.4]
  input  [31:0] io_input_regs_2_a4, // @[:@6.4]
  input  [31:0] io_input_regs_2_a5, // @[:@6.4]
  input  [31:0] io_input_regs_2_a6, // @[:@6.4]
  input  [31:0] io_input_regs_2_a7, // @[:@6.4]
  input  [31:0] io_input_regs_2_s2, // @[:@6.4]
  input  [31:0] io_input_regs_2_s3, // @[:@6.4]
  input  [31:0] io_input_regs_2_s4, // @[:@6.4]
  input  [31:0] io_input_regs_2_s5, // @[:@6.4]
  input  [31:0] io_input_regs_2_s6, // @[:@6.4]
  input  [31:0] io_input_regs_2_s7, // @[:@6.4]
  input  [31:0] io_input_regs_2_s8, // @[:@6.4]
  input  [31:0] io_input_regs_2_s9, // @[:@6.4]
  input  [31:0] io_input_regs_2_s10, // @[:@6.4]
  input  [31:0] io_input_regs_2_s11, // @[:@6.4]
  input  [31:0] io_input_regs_2_t3, // @[:@6.4]
  input  [31:0] io_input_regs_2_t4, // @[:@6.4]
  input  [31:0] io_input_regs_2_t5, // @[:@6.4]
  input  [31:0] io_input_regs_2_t6, // @[:@6.4]
  input  [31:0] io_input_regs_2_pc, // @[:@6.4]
  input         io_input_regs_2_interrupt, // @[:@6.4]
  input  [31:0] io_input_regs_2_interrupt_cause, // @[:@6.4]
  input  [31:0] io_input_regs_2_time, // @[:@6.4]
  input         io_input_regs_2_debug, // @[:@6.4]
  input  [31:0] io_input_regs_2_isa, // @[:@6.4]
  input         io_input_regs_2_sd, // @[:@6.4]
  input         io_input_regs_2_sd_rv32, // @[:@6.4]
  input  [31:0] io_input_regs_2_mpp, // @[:@6.4]
  input         io_input_regs_2_spp, // @[:@6.4]
  input         io_input_regs_2_mpie, // @[:@6.4]
  input         io_input_regs_2_mie, // @[:@6.4]
  input  [31:0] io_input_regs_2_evec, // @[:@6.4]
  output [31:0] io_output_regs_0_ra, // @[:@6.4]
  output [31:0] io_output_regs_0_sp, // @[:@6.4]
  output [31:0] io_output_regs_0_gp, // @[:@6.4]
  output [31:0] io_output_regs_0_tp, // @[:@6.4]
  output [31:0] io_output_regs_0_t0, // @[:@6.4]
  output [31:0] io_output_regs_0_t1, // @[:@6.4]
  output [31:0] io_output_regs_0_t2, // @[:@6.4]
  output [31:0] io_output_regs_0_fp, // @[:@6.4]
  output [31:0] io_output_regs_0_s1, // @[:@6.4]
  output [31:0] io_output_regs_0_a0, // @[:@6.4]
  output [31:0] io_output_regs_0_a1, // @[:@6.4]
  output [31:0] io_output_regs_0_a2, // @[:@6.4]
  output [31:0] io_output_regs_0_a3, // @[:@6.4]
  output [31:0] io_output_regs_0_a4, // @[:@6.4]
  output [31:0] io_output_regs_0_a5, // @[:@6.4]
  output [31:0] io_output_regs_0_a6, // @[:@6.4]
  output [31:0] io_output_regs_0_a7, // @[:@6.4]
  output [31:0] io_output_regs_0_s2, // @[:@6.4]
  output [31:0] io_output_regs_0_s3, // @[:@6.4]
  output [31:0] io_output_regs_0_s4, // @[:@6.4]
  output [31:0] io_output_regs_0_s5, // @[:@6.4]
  output [31:0] io_output_regs_0_s6, // @[:@6.4]
  output [31:0] io_output_regs_0_s7, // @[:@6.4]
  output [31:0] io_output_regs_0_s8, // @[:@6.4]
  output [31:0] io_output_regs_0_s9, // @[:@6.4]
  output [31:0] io_output_regs_0_s10, // @[:@6.4]
  output [31:0] io_output_regs_0_s11, // @[:@6.4]
  output [31:0] io_output_regs_0_t3, // @[:@6.4]
  output [31:0] io_output_regs_0_t4, // @[:@6.4]
  output [31:0] io_output_regs_0_t5, // @[:@6.4]
  output [31:0] io_output_regs_0_t6, // @[:@6.4]
  output [31:0] io_output_regs_0_pc, // @[:@6.4]
  output        io_output_regs_0_interrupt, // @[:@6.4]
  output [31:0] io_output_regs_0_interrupt_cause, // @[:@6.4]
  output [31:0] io_output_regs_0_time, // @[:@6.4]
  output        io_output_regs_0_debug, // @[:@6.4]
  output [31:0] io_output_regs_0_isa, // @[:@6.4]
  output        io_output_regs_0_sd, // @[:@6.4]
  output        io_output_regs_0_sd_rv32, // @[:@6.4]
  output [31:0] io_output_regs_0_mpp, // @[:@6.4]
  output        io_output_regs_0_spp, // @[:@6.4]
  output        io_output_regs_0_mpie, // @[:@6.4]
  output        io_output_regs_0_mie, // @[:@6.4]
  output [31:0] io_output_regs_0_evec, // @[:@6.4]
  output [31:0] io_output_regs_1_ra, // @[:@6.4]
  output [31:0] io_output_regs_1_sp, // @[:@6.4]
  output [31:0] io_output_regs_1_gp, // @[:@6.4]
  output [31:0] io_output_regs_1_tp, // @[:@6.4]
  output [31:0] io_output_regs_1_t0, // @[:@6.4]
  output [31:0] io_output_regs_1_t1, // @[:@6.4]
  output [31:0] io_output_regs_1_t2, // @[:@6.4]
  output [31:0] io_output_regs_1_fp, // @[:@6.4]
  output [31:0] io_output_regs_1_s1, // @[:@6.4]
  output [31:0] io_output_regs_1_a0, // @[:@6.4]
  output [31:0] io_output_regs_1_a1, // @[:@6.4]
  output [31:0] io_output_regs_1_a2, // @[:@6.4]
  output [31:0] io_output_regs_1_a3, // @[:@6.4]
  output [31:0] io_output_regs_1_a4, // @[:@6.4]
  output [31:0] io_output_regs_1_a5, // @[:@6.4]
  output [31:0] io_output_regs_1_a6, // @[:@6.4]
  output [31:0] io_output_regs_1_a7, // @[:@6.4]
  output [31:0] io_output_regs_1_s2, // @[:@6.4]
  output [31:0] io_output_regs_1_s3, // @[:@6.4]
  output [31:0] io_output_regs_1_s4, // @[:@6.4]
  output [31:0] io_output_regs_1_s5, // @[:@6.4]
  output [31:0] io_output_regs_1_s6, // @[:@6.4]
  output [31:0] io_output_regs_1_s7, // @[:@6.4]
  output [31:0] io_output_regs_1_s8, // @[:@6.4]
  output [31:0] io_output_regs_1_s9, // @[:@6.4]
  output [31:0] io_output_regs_1_s10, // @[:@6.4]
  output [31:0] io_output_regs_1_s11, // @[:@6.4]
  output [31:0] io_output_regs_1_t3, // @[:@6.4]
  output [31:0] io_output_regs_1_t4, // @[:@6.4]
  output [31:0] io_output_regs_1_t5, // @[:@6.4]
  output [31:0] io_output_regs_1_t6, // @[:@6.4]
  output [31:0] io_output_regs_1_pc, // @[:@6.4]
  output        io_output_regs_1_interrupt, // @[:@6.4]
  output [31:0] io_output_regs_1_interrupt_cause, // @[:@6.4]
  output [31:0] io_output_regs_1_time, // @[:@6.4]
  output        io_output_regs_1_debug, // @[:@6.4]
  output [31:0] io_output_regs_1_isa, // @[:@6.4]
  output        io_output_regs_1_sd, // @[:@6.4]
  output        io_output_regs_1_sd_rv32, // @[:@6.4]
  output [31:0] io_output_regs_1_mpp, // @[:@6.4]
  output        io_output_regs_1_spp, // @[:@6.4]
  output        io_output_regs_1_mpie, // @[:@6.4]
  output        io_output_regs_1_mie, // @[:@6.4]
  output [31:0] io_output_regs_1_evec, // @[:@6.4]
  output [31:0] io_output_regs_2_ra, // @[:@6.4]
  output [31:0] io_output_regs_2_sp, // @[:@6.4]
  output [31:0] io_output_regs_2_gp, // @[:@6.4]
  output [31:0] io_output_regs_2_tp, // @[:@6.4]
  output [31:0] io_output_regs_2_t0, // @[:@6.4]
  output [31:0] io_output_regs_2_t1, // @[:@6.4]
  output [31:0] io_output_regs_2_t2, // @[:@6.4]
  output [31:0] io_output_regs_2_fp, // @[:@6.4]
  output [31:0] io_output_regs_2_s1, // @[:@6.4]
  output [31:0] io_output_regs_2_a0, // @[:@6.4]
  output [31:0] io_output_regs_2_a1, // @[:@6.4]
  output [31:0] io_output_regs_2_a2, // @[:@6.4]
  output [31:0] io_output_regs_2_a3, // @[:@6.4]
  output [31:0] io_output_regs_2_a4, // @[:@6.4]
  output [31:0] io_output_regs_2_a5, // @[:@6.4]
  output [31:0] io_output_regs_2_a6, // @[:@6.4]
  output [31:0] io_output_regs_2_a7, // @[:@6.4]
  output [31:0] io_output_regs_2_s2, // @[:@6.4]
  output [31:0] io_output_regs_2_s3, // @[:@6.4]
  output [31:0] io_output_regs_2_s4, // @[:@6.4]
  output [31:0] io_output_regs_2_s5, // @[:@6.4]
  output [31:0] io_output_regs_2_s6, // @[:@6.4]
  output [31:0] io_output_regs_2_s7, // @[:@6.4]
  output [31:0] io_output_regs_2_s8, // @[:@6.4]
  output [31:0] io_output_regs_2_s9, // @[:@6.4]
  output [31:0] io_output_regs_2_s10, // @[:@6.4]
  output [31:0] io_output_regs_2_s11, // @[:@6.4]
  output [31:0] io_output_regs_2_t3, // @[:@6.4]
  output [31:0] io_output_regs_2_t4, // @[:@6.4]
  output [31:0] io_output_regs_2_t5, // @[:@6.4]
  output [31:0] io_output_regs_2_t6, // @[:@6.4]
  output [31:0] io_output_regs_2_pc, // @[:@6.4]
  output        io_output_regs_2_interrupt, // @[:@6.4]
  output [31:0] io_output_regs_2_interrupt_cause, // @[:@6.4]
  output [31:0] io_output_regs_2_time, // @[:@6.4]
  output        io_output_regs_2_debug, // @[:@6.4]
  output [31:0] io_output_regs_2_isa, // @[:@6.4]
  output        io_output_regs_2_sd, // @[:@6.4]
  output        io_output_regs_2_sd_rv32, // @[:@6.4]
  output [31:0] io_output_regs_2_mpp, // @[:@6.4]
  output        io_output_regs_2_spp, // @[:@6.4]
  output        io_output_regs_2_mpie, // @[:@6.4]
  output        io_output_regs_2_mie, // @[:@6.4]
  output [31:0] io_output_regs_2_evec // @[:@6.4]
);
  wire  _T_985; // @[RegsRouter.scala 68:20:@8.4]
  wire [31:0] _T_986; // @[RegsRouter.scala 10:33:@10.6]
  wire [31:0] _T_987; // @[RegsRouter.scala 11:33:@12.6]
  wire [31:0] _T_988; // @[RegsRouter.scala 12:33:@14.6]
  wire [31:0] _T_989; // @[RegsRouter.scala 13:33:@16.6]
  wire [31:0] _T_990; // @[RegsRouter.scala 14:33:@18.6]
  wire [31:0] _T_991; // @[RegsRouter.scala 15:33:@20.6]
  wire [31:0] _T_992; // @[RegsRouter.scala 16:33:@22.6]
  wire [31:0] _T_993; // @[RegsRouter.scala 17:33:@24.6]
  wire [31:0] _T_994; // @[RegsRouter.scala 18:33:@26.6]
  wire [31:0] _T_995; // @[RegsRouter.scala 19:33:@28.6]
  wire [31:0] _T_996; // @[RegsRouter.scala 20:33:@30.6]
  wire [31:0] _T_997; // @[RegsRouter.scala 21:33:@32.6]
  wire [31:0] _T_998; // @[RegsRouter.scala 22:33:@34.6]
  wire [31:0] _T_999; // @[RegsRouter.scala 23:33:@36.6]
  wire [31:0] _T_1000; // @[RegsRouter.scala 24:33:@38.6]
  wire [31:0] _T_1001; // @[RegsRouter.scala 25:33:@40.6]
  wire [31:0] _T_1002; // @[RegsRouter.scala 26:33:@42.6]
  wire [31:0] _T_1003; // @[RegsRouter.scala 27:33:@44.6]
  wire [31:0] _T_1004; // @[RegsRouter.scala 28:33:@46.6]
  wire [31:0] _T_1005; // @[RegsRouter.scala 29:33:@48.6]
  wire [31:0] _T_1006; // @[RegsRouter.scala 30:33:@50.6]
  wire [31:0] _T_1007; // @[RegsRouter.scala 31:33:@52.6]
  wire [31:0] _T_1008; // @[RegsRouter.scala 32:33:@54.6]
  wire [31:0] _T_1009; // @[RegsRouter.scala 33:33:@56.6]
  wire [31:0] _T_1010; // @[RegsRouter.scala 34:33:@58.6]
  wire [31:0] _T_1011; // @[RegsRouter.scala 35:35:@60.6]
  wire [31:0] _T_1012; // @[RegsRouter.scala 36:35:@62.6]
  wire [31:0] _T_1013; // @[RegsRouter.scala 37:33:@64.6]
  wire [31:0] _T_1014; // @[RegsRouter.scala 38:33:@66.6]
  wire [31:0] _T_1015; // @[RegsRouter.scala 39:33:@68.6]
  wire [31:0] _T_1016; // @[RegsRouter.scala 40:33:@70.6]
  wire [31:0] _T_1017; // @[RegsRouter.scala 41:33:@72.6]
  wire  _T_1018; // @[RegsRouter.scala 42:47:@74.6]
  wire [31:0] _T_1019; // @[RegsRouter.scala 43:59:@76.6]
  wire [31:0] _T_1020; // @[RegsRouter.scala 44:37:@78.6]
  wire  _T_1021; // @[RegsRouter.scala 45:39:@80.6]
  wire [31:0] _T_1022; // @[RegsRouter.scala 46:35:@82.6]
  wire  _T_1023; // @[RegsRouter.scala 47:33:@84.6]
  wire  _T_1024; // @[RegsRouter.scala 48:43:@86.6]
  wire [31:0] _T_1025; // @[RegsRouter.scala 49:35:@88.6]
  wire  _T_1026; // @[RegsRouter.scala 50:35:@90.6]
  wire  _T_1027; // @[RegsRouter.scala 51:37:@92.6]
  wire  _T_1028; // @[RegsRouter.scala 52:35:@94.6]
  wire [31:0] _T_1029; // @[RegsRouter.scala 53:37:@96.6]
  wire [31:0] _T_1030; // @[RegsRouter.scala 10:33:@98.6]
  wire [31:0] _T_1031; // @[RegsRouter.scala 11:33:@100.6]
  wire [31:0] _T_1032; // @[RegsRouter.scala 12:33:@102.6]
  wire [31:0] _T_1033; // @[RegsRouter.scala 13:33:@104.6]
  wire [31:0] _T_1034; // @[RegsRouter.scala 14:33:@106.6]
  wire [31:0] _T_1035; // @[RegsRouter.scala 15:33:@108.6]
  wire [31:0] _T_1036; // @[RegsRouter.scala 16:33:@110.6]
  wire [31:0] _T_1037; // @[RegsRouter.scala 17:33:@112.6]
  wire [31:0] _T_1038; // @[RegsRouter.scala 18:33:@114.6]
  wire [31:0] _T_1039; // @[RegsRouter.scala 19:33:@116.6]
  wire [31:0] _T_1040; // @[RegsRouter.scala 20:33:@118.6]
  wire [31:0] _T_1041; // @[RegsRouter.scala 21:33:@120.6]
  wire [31:0] _T_1042; // @[RegsRouter.scala 22:33:@122.6]
  wire [31:0] _T_1043; // @[RegsRouter.scala 23:33:@124.6]
  wire [31:0] _T_1044; // @[RegsRouter.scala 24:33:@126.6]
  wire [31:0] _T_1045; // @[RegsRouter.scala 25:33:@128.6]
  wire [31:0] _T_1046; // @[RegsRouter.scala 26:33:@130.6]
  wire [31:0] _T_1047; // @[RegsRouter.scala 27:33:@132.6]
  wire [31:0] _T_1048; // @[RegsRouter.scala 28:33:@134.6]
  wire [31:0] _T_1049; // @[RegsRouter.scala 29:33:@136.6]
  wire [31:0] _T_1050; // @[RegsRouter.scala 30:33:@138.6]
  wire [31:0] _T_1051; // @[RegsRouter.scala 31:33:@140.6]
  wire [31:0] _T_1052; // @[RegsRouter.scala 32:33:@142.6]
  wire [31:0] _T_1053; // @[RegsRouter.scala 33:33:@144.6]
  wire [31:0] _T_1054; // @[RegsRouter.scala 34:33:@146.6]
  wire [31:0] _T_1055; // @[RegsRouter.scala 35:35:@148.6]
  wire [31:0] _T_1056; // @[RegsRouter.scala 36:35:@150.6]
  wire [31:0] _T_1057; // @[RegsRouter.scala 37:33:@152.6]
  wire [31:0] _T_1058; // @[RegsRouter.scala 38:33:@154.6]
  wire [31:0] _T_1059; // @[RegsRouter.scala 39:33:@156.6]
  wire [31:0] _T_1060; // @[RegsRouter.scala 40:33:@158.6]
  wire [31:0] _T_1061; // @[RegsRouter.scala 41:33:@160.6]
  wire  _T_1062; // @[RegsRouter.scala 42:47:@162.6]
  wire [31:0] _T_1063; // @[RegsRouter.scala 43:59:@164.6]
  wire [31:0] _T_1064; // @[RegsRouter.scala 44:37:@166.6]
  wire  _T_1065; // @[RegsRouter.scala 45:39:@168.6]
  wire [31:0] _T_1066; // @[RegsRouter.scala 46:35:@170.6]
  wire  _T_1067; // @[RegsRouter.scala 47:33:@172.6]
  wire  _T_1068; // @[RegsRouter.scala 48:43:@174.6]
  wire [31:0] _T_1069; // @[RegsRouter.scala 49:35:@176.6]
  wire  _T_1070; // @[RegsRouter.scala 50:35:@178.6]
  wire  _T_1071; // @[RegsRouter.scala 51:37:@180.6]
  wire  _T_1072; // @[RegsRouter.scala 52:35:@182.6]
  wire [31:0] _T_1073; // @[RegsRouter.scala 53:37:@184.6]
  wire [31:0] _T_1074; // @[RegsRouter.scala 10:33:@186.6]
  wire [31:0] _T_1075; // @[RegsRouter.scala 11:33:@188.6]
  wire [31:0] _T_1076; // @[RegsRouter.scala 12:33:@190.6]
  wire [31:0] _T_1077; // @[RegsRouter.scala 13:33:@192.6]
  wire [31:0] _T_1078; // @[RegsRouter.scala 14:33:@194.6]
  wire [31:0] _T_1079; // @[RegsRouter.scala 15:33:@196.6]
  wire [31:0] _T_1080; // @[RegsRouter.scala 16:33:@198.6]
  wire [31:0] _T_1081; // @[RegsRouter.scala 17:33:@200.6]
  wire [31:0] _T_1082; // @[RegsRouter.scala 18:33:@202.6]
  wire [31:0] _T_1083; // @[RegsRouter.scala 19:33:@204.6]
  wire [31:0] _T_1084; // @[RegsRouter.scala 20:33:@206.6]
  wire [31:0] _T_1085; // @[RegsRouter.scala 21:33:@208.6]
  wire [31:0] _T_1086; // @[RegsRouter.scala 22:33:@210.6]
  wire [31:0] _T_1087; // @[RegsRouter.scala 23:33:@212.6]
  wire [31:0] _T_1088; // @[RegsRouter.scala 24:33:@214.6]
  wire [31:0] _T_1089; // @[RegsRouter.scala 25:33:@216.6]
  wire [31:0] _T_1090; // @[RegsRouter.scala 26:33:@218.6]
  wire [31:0] _T_1091; // @[RegsRouter.scala 27:33:@220.6]
  wire [31:0] _T_1092; // @[RegsRouter.scala 28:33:@222.6]
  wire [31:0] _T_1093; // @[RegsRouter.scala 29:33:@224.6]
  wire [31:0] _T_1094; // @[RegsRouter.scala 30:33:@226.6]
  wire [31:0] _T_1095; // @[RegsRouter.scala 31:33:@228.6]
  wire [31:0] _T_1096; // @[RegsRouter.scala 32:33:@230.6]
  wire [31:0] _T_1097; // @[RegsRouter.scala 33:33:@232.6]
  wire [31:0] _T_1098; // @[RegsRouter.scala 34:33:@234.6]
  wire [31:0] _T_1099; // @[RegsRouter.scala 35:35:@236.6]
  wire [31:0] _T_1100; // @[RegsRouter.scala 36:35:@238.6]
  wire [31:0] _T_1101; // @[RegsRouter.scala 37:33:@240.6]
  wire [31:0] _T_1102; // @[RegsRouter.scala 38:33:@242.6]
  wire [31:0] _T_1103; // @[RegsRouter.scala 39:33:@244.6]
  wire [31:0] _T_1104; // @[RegsRouter.scala 40:33:@246.6]
  wire [31:0] _T_1105; // @[RegsRouter.scala 41:33:@248.6]
  wire  _T_1106; // @[RegsRouter.scala 42:47:@250.6]
  wire [31:0] _T_1107; // @[RegsRouter.scala 43:59:@252.6]
  wire [31:0] _T_1108; // @[RegsRouter.scala 44:37:@254.6]
  wire  _T_1109; // @[RegsRouter.scala 45:39:@256.6]
  wire [31:0] _T_1110; // @[RegsRouter.scala 46:35:@258.6]
  wire  _T_1111; // @[RegsRouter.scala 47:33:@260.6]
  wire  _T_1112; // @[RegsRouter.scala 48:43:@262.6]
  wire [31:0] _T_1113; // @[RegsRouter.scala 49:35:@264.6]
  wire  _T_1114; // @[RegsRouter.scala 50:35:@266.6]
  wire  _T_1115; // @[RegsRouter.scala 51:37:@268.6]
  wire  _T_1116; // @[RegsRouter.scala 52:35:@270.6]
  wire [31:0] _T_1117; // @[RegsRouter.scala 53:37:@272.6]
  wire  _T_1118; // @[RegsRouter.scala 73:26:@276.6]
  wire [31:0] _T_1119; // @[RegsRouter.scala 10:33:@278.8]
  wire [31:0] _T_1120; // @[RegsRouter.scala 11:33:@280.8]
  wire [31:0] _T_1121; // @[RegsRouter.scala 12:33:@282.8]
  wire [31:0] _T_1122; // @[RegsRouter.scala 13:33:@284.8]
  wire [31:0] _T_1123; // @[RegsRouter.scala 14:33:@286.8]
  wire [31:0] _T_1124; // @[RegsRouter.scala 15:33:@288.8]
  wire [31:0] _T_1125; // @[RegsRouter.scala 16:33:@290.8]
  wire [31:0] _T_1126; // @[RegsRouter.scala 17:33:@292.8]
  wire [31:0] _T_1127; // @[RegsRouter.scala 18:33:@294.8]
  wire [31:0] _T_1128; // @[RegsRouter.scala 19:33:@296.8]
  wire [31:0] _T_1129; // @[RegsRouter.scala 20:33:@298.8]
  wire [31:0] _T_1130; // @[RegsRouter.scala 21:33:@300.8]
  wire [31:0] _T_1131; // @[RegsRouter.scala 22:33:@302.8]
  wire [31:0] _T_1132; // @[RegsRouter.scala 23:33:@304.8]
  wire [31:0] _T_1133; // @[RegsRouter.scala 24:33:@306.8]
  wire [31:0] _T_1134; // @[RegsRouter.scala 25:33:@308.8]
  wire [31:0] _T_1135; // @[RegsRouter.scala 26:33:@310.8]
  wire [31:0] _T_1136; // @[RegsRouter.scala 27:33:@312.8]
  wire [31:0] _T_1137; // @[RegsRouter.scala 28:33:@314.8]
  wire [31:0] _T_1138; // @[RegsRouter.scala 29:33:@316.8]
  wire [31:0] _T_1139; // @[RegsRouter.scala 30:33:@318.8]
  wire [31:0] _T_1140; // @[RegsRouter.scala 31:33:@320.8]
  wire [31:0] _T_1141; // @[RegsRouter.scala 32:33:@322.8]
  wire [31:0] _T_1142; // @[RegsRouter.scala 33:33:@324.8]
  wire [31:0] _T_1143; // @[RegsRouter.scala 34:33:@326.8]
  wire [31:0] _T_1144; // @[RegsRouter.scala 35:35:@328.8]
  wire [31:0] _T_1145; // @[RegsRouter.scala 36:35:@330.8]
  wire [31:0] _T_1146; // @[RegsRouter.scala 37:33:@332.8]
  wire [31:0] _T_1147; // @[RegsRouter.scala 38:33:@334.8]
  wire [31:0] _T_1148; // @[RegsRouter.scala 39:33:@336.8]
  wire [31:0] _T_1149; // @[RegsRouter.scala 40:33:@338.8]
  wire [31:0] _T_1150; // @[RegsRouter.scala 41:33:@340.8]
  wire  _T_1151; // @[RegsRouter.scala 42:47:@342.8]
  wire [31:0] _T_1152; // @[RegsRouter.scala 43:59:@344.8]
  wire [31:0] _T_1153; // @[RegsRouter.scala 44:37:@346.8]
  wire  _T_1154; // @[RegsRouter.scala 45:39:@348.8]
  wire [31:0] _T_1155; // @[RegsRouter.scala 46:35:@350.8]
  wire  _T_1156; // @[RegsRouter.scala 47:33:@352.8]
  wire  _T_1157; // @[RegsRouter.scala 48:43:@354.8]
  wire [31:0] _T_1158; // @[RegsRouter.scala 49:35:@356.8]
  wire  _T_1159; // @[RegsRouter.scala 50:35:@358.8]
  wire  _T_1160; // @[RegsRouter.scala 51:37:@360.8]
  wire  _T_1161; // @[RegsRouter.scala 52:35:@362.8]
  wire [31:0] _T_1162; // @[RegsRouter.scala 53:37:@364.8]
  wire [31:0] _T_1163; // @[RegsRouter.scala 10:33:@366.8]
  wire [31:0] _T_1164; // @[RegsRouter.scala 11:33:@368.8]
  wire [31:0] _T_1165; // @[RegsRouter.scala 12:33:@370.8]
  wire [31:0] _T_1166; // @[RegsRouter.scala 13:33:@372.8]
  wire [31:0] _T_1167; // @[RegsRouter.scala 14:33:@374.8]
  wire [31:0] _T_1168; // @[RegsRouter.scala 15:33:@376.8]
  wire [31:0] _T_1169; // @[RegsRouter.scala 16:33:@378.8]
  wire [31:0] _T_1170; // @[RegsRouter.scala 17:33:@380.8]
  wire [31:0] _T_1171; // @[RegsRouter.scala 18:33:@382.8]
  wire [31:0] _T_1172; // @[RegsRouter.scala 19:33:@384.8]
  wire [31:0] _T_1173; // @[RegsRouter.scala 20:33:@386.8]
  wire [31:0] _T_1174; // @[RegsRouter.scala 21:33:@388.8]
  wire [31:0] _T_1175; // @[RegsRouter.scala 22:33:@390.8]
  wire [31:0] _T_1176; // @[RegsRouter.scala 23:33:@392.8]
  wire [31:0] _T_1177; // @[RegsRouter.scala 24:33:@394.8]
  wire [31:0] _T_1178; // @[RegsRouter.scala 25:33:@396.8]
  wire [31:0] _T_1179; // @[RegsRouter.scala 26:33:@398.8]
  wire [31:0] _T_1180; // @[RegsRouter.scala 27:33:@400.8]
  wire [31:0] _T_1181; // @[RegsRouter.scala 28:33:@402.8]
  wire [31:0] _T_1182; // @[RegsRouter.scala 29:33:@404.8]
  wire [31:0] _T_1183; // @[RegsRouter.scala 30:33:@406.8]
  wire [31:0] _T_1184; // @[RegsRouter.scala 31:33:@408.8]
  wire [31:0] _T_1185; // @[RegsRouter.scala 32:33:@410.8]
  wire [31:0] _T_1186; // @[RegsRouter.scala 33:33:@412.8]
  wire [31:0] _T_1187; // @[RegsRouter.scala 34:33:@414.8]
  wire [31:0] _T_1188; // @[RegsRouter.scala 35:35:@416.8]
  wire [31:0] _T_1189; // @[RegsRouter.scala 36:35:@418.8]
  wire [31:0] _T_1190; // @[RegsRouter.scala 37:33:@420.8]
  wire [31:0] _T_1191; // @[RegsRouter.scala 38:33:@422.8]
  wire [31:0] _T_1192; // @[RegsRouter.scala 39:33:@424.8]
  wire [31:0] _T_1193; // @[RegsRouter.scala 40:33:@426.8]
  wire [31:0] _T_1194; // @[RegsRouter.scala 41:33:@428.8]
  wire  _T_1195; // @[RegsRouter.scala 42:47:@430.8]
  wire [31:0] _T_1196; // @[RegsRouter.scala 43:59:@432.8]
  wire [31:0] _T_1197; // @[RegsRouter.scala 44:37:@434.8]
  wire  _T_1198; // @[RegsRouter.scala 45:39:@436.8]
  wire [31:0] _T_1199; // @[RegsRouter.scala 46:35:@438.8]
  wire  _T_1200; // @[RegsRouter.scala 47:33:@440.8]
  wire  _T_1201; // @[RegsRouter.scala 48:43:@442.8]
  wire [31:0] _T_1202; // @[RegsRouter.scala 49:35:@444.8]
  wire  _T_1203; // @[RegsRouter.scala 50:35:@446.8]
  wire  _T_1204; // @[RegsRouter.scala 51:37:@448.8]
  wire  _T_1205; // @[RegsRouter.scala 52:35:@450.8]
  wire [31:0] _T_1206; // @[RegsRouter.scala 53:37:@452.8]
  wire  _T_1251; // @[RegsRouter.scala 78:26:@544.8]
  wire [31:0] _T_1340; // @[RegsRouter.scala 10:33:@722.10]
  wire [31:0] _T_1341; // @[RegsRouter.scala 11:33:@724.10]
  wire [31:0] _T_1342; // @[RegsRouter.scala 12:33:@726.10]
  wire [31:0] _T_1343; // @[RegsRouter.scala 13:33:@728.10]
  wire [31:0] _T_1344; // @[RegsRouter.scala 14:33:@730.10]
  wire [31:0] _T_1345; // @[RegsRouter.scala 15:33:@732.10]
  wire [31:0] _T_1346; // @[RegsRouter.scala 16:33:@734.10]
  wire [31:0] _T_1347; // @[RegsRouter.scala 17:33:@736.10]
  wire [31:0] _T_1348; // @[RegsRouter.scala 18:33:@738.10]
  wire [31:0] _T_1349; // @[RegsRouter.scala 19:33:@740.10]
  wire [31:0] _T_1350; // @[RegsRouter.scala 20:33:@742.10]
  wire [31:0] _T_1351; // @[RegsRouter.scala 21:33:@744.10]
  wire [31:0] _T_1352; // @[RegsRouter.scala 22:33:@746.10]
  wire [31:0] _T_1353; // @[RegsRouter.scala 23:33:@748.10]
  wire [31:0] _T_1354; // @[RegsRouter.scala 24:33:@750.10]
  wire [31:0] _T_1355; // @[RegsRouter.scala 25:33:@752.10]
  wire [31:0] _T_1356; // @[RegsRouter.scala 26:33:@754.10]
  wire [31:0] _T_1357; // @[RegsRouter.scala 27:33:@756.10]
  wire [31:0] _T_1358; // @[RegsRouter.scala 28:33:@758.10]
  wire [31:0] _T_1359; // @[RegsRouter.scala 29:33:@760.10]
  wire [31:0] _T_1360; // @[RegsRouter.scala 30:33:@762.10]
  wire [31:0] _T_1361; // @[RegsRouter.scala 31:33:@764.10]
  wire [31:0] _T_1362; // @[RegsRouter.scala 32:33:@766.10]
  wire [31:0] _T_1363; // @[RegsRouter.scala 33:33:@768.10]
  wire [31:0] _T_1364; // @[RegsRouter.scala 34:33:@770.10]
  wire [31:0] _T_1365; // @[RegsRouter.scala 35:35:@772.10]
  wire [31:0] _T_1366; // @[RegsRouter.scala 36:35:@774.10]
  wire [31:0] _T_1367; // @[RegsRouter.scala 37:33:@776.10]
  wire [31:0] _T_1368; // @[RegsRouter.scala 38:33:@778.10]
  wire [31:0] _T_1369; // @[RegsRouter.scala 39:33:@780.10]
  wire [31:0] _T_1370; // @[RegsRouter.scala 40:33:@782.10]
  wire [31:0] _T_1371; // @[RegsRouter.scala 41:33:@784.10]
  wire  _T_1372; // @[RegsRouter.scala 42:47:@786.10]
  wire [31:0] _T_1373; // @[RegsRouter.scala 43:59:@788.10]
  wire [31:0] _T_1374; // @[RegsRouter.scala 44:37:@790.10]
  wire  _T_1375; // @[RegsRouter.scala 45:39:@792.10]
  wire [31:0] _T_1376; // @[RegsRouter.scala 46:35:@794.10]
  wire  _T_1377; // @[RegsRouter.scala 47:33:@796.10]
  wire  _T_1378; // @[RegsRouter.scala 48:43:@798.10]
  wire [31:0] _T_1379; // @[RegsRouter.scala 49:35:@800.10]
  wire  _T_1380; // @[RegsRouter.scala 50:35:@802.10]
  wire  _T_1381; // @[RegsRouter.scala 51:37:@804.10]
  wire  _T_1382; // @[RegsRouter.scala 52:35:@806.10]
  wire [31:0] _T_1383; // @[RegsRouter.scala 53:37:@808.10]
  wire [31:0] _GEN_0; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_1; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_2; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_3; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_4; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_5; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_6; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_7; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_8; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_9; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_10; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_11; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_12; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_13; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_14; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_15; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_16; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_17; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_18; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_19; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_20; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_21; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_22; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_23; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_24; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_25; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_26; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_27; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_28; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_29; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_30; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_31; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_32; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_33; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_34; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_35; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_36; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_37; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_38; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_39; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_40; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_41; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_42; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_43; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_44; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_45; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_46; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_47; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_48; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_49; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_50; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_51; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_52; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_53; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_54; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_55; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_56; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_57; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_58; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_59; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_60; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_61; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_62; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_63; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_64; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_65; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_66; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_67; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_68; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_69; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_70; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_71; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_72; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_73; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_74; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_75; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_76; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_77; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_78; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_79; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_80; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_81; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_82; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_83; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_84; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_85; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_86; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_87; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_88; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_89; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_90; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_91; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_92; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_93; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_94; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_95; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_96; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_97; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_98; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_99; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_100; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_101; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_102; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_103; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_104; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_105; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_106; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_107; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_108; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_109; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_110; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_111; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_112; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_113; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_114; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_115; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_116; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_117; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_118; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_119; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_120; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_121; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_122; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_123; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_124; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_125; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_126; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_127; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_128; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_129; // @[RegsRouter.scala 78:44:@545.8]
  wire  _GEN_130; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_131; // @[RegsRouter.scala 78:44:@545.8]
  wire [31:0] _GEN_132; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_133; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_134; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_135; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_136; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_137; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_138; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_139; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_140; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_141; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_142; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_143; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_144; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_145; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_146; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_147; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_148; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_149; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_150; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_151; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_152; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_153; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_154; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_155; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_156; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_157; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_158; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_159; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_160; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_161; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_162; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_163; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_164; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_165; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_166; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_167; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_168; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_169; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_170; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_171; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_172; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_173; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_174; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_175; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_176; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_177; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_178; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_179; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_180; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_181; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_182; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_183; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_184; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_185; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_186; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_187; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_188; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_189; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_190; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_191; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_192; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_193; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_194; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_195; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_196; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_197; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_198; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_199; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_200; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_201; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_202; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_203; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_204; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_205; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_206; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_207; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_208; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_209; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_210; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_211; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_212; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_213; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_214; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_215; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_216; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_217; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_218; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_219; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_220; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_221; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_222; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_223; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_224; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_225; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_226; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_227; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_228; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_229; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_230; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_231; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_232; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_233; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_234; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_235; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_236; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_237; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_238; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_239; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_240; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_241; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_242; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_243; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_244; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_245; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_246; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_247; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_248; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_249; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_250; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_251; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_252; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_253; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_254; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_255; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_256; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_257; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_258; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_259; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_260; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_261; // @[RegsRouter.scala 73:44:@277.6]
  wire  _GEN_262; // @[RegsRouter.scala 73:44:@277.6]
  wire [31:0] _GEN_263; // @[RegsRouter.scala 73:44:@277.6]
  assign _T_985 = io_selector == 3'h1; // @[RegsRouter.scala 68:20:@8.4]
  assign _T_986 = io_input_regs_1_ra | io_input_regs_2_ra; // @[RegsRouter.scala 10:33:@10.6]
  assign _T_987 = io_input_regs_1_sp | io_input_regs_2_sp; // @[RegsRouter.scala 11:33:@12.6]
  assign _T_988 = io_input_regs_1_gp | io_input_regs_2_gp; // @[RegsRouter.scala 12:33:@14.6]
  assign _T_989 = io_input_regs_1_tp | io_input_regs_2_tp; // @[RegsRouter.scala 13:33:@16.6]
  assign _T_990 = io_input_regs_1_t0 | io_input_regs_2_t0; // @[RegsRouter.scala 14:33:@18.6]
  assign _T_991 = io_input_regs_1_t1 | io_input_regs_2_t1; // @[RegsRouter.scala 15:33:@20.6]
  assign _T_992 = io_input_regs_1_t2 | io_input_regs_2_t2; // @[RegsRouter.scala 16:33:@22.6]
  assign _T_993 = io_input_regs_1_fp | io_input_regs_2_fp; // @[RegsRouter.scala 17:33:@24.6]
  assign _T_994 = io_input_regs_1_s1 | io_input_regs_2_s1; // @[RegsRouter.scala 18:33:@26.6]
  assign _T_995 = io_input_regs_1_a0 | io_input_regs_2_a0; // @[RegsRouter.scala 19:33:@28.6]
  assign _T_996 = io_input_regs_1_a1 | io_input_regs_2_a1; // @[RegsRouter.scala 20:33:@30.6]
  assign _T_997 = io_input_regs_1_a2 | io_input_regs_2_a2; // @[RegsRouter.scala 21:33:@32.6]
  assign _T_998 = io_input_regs_1_a3 | io_input_regs_2_a3; // @[RegsRouter.scala 22:33:@34.6]
  assign _T_999 = io_input_regs_1_a4 | io_input_regs_2_a4; // @[RegsRouter.scala 23:33:@36.6]
  assign _T_1000 = io_input_regs_1_a5 | io_input_regs_2_a5; // @[RegsRouter.scala 24:33:@38.6]
  assign _T_1001 = io_input_regs_1_a6 | io_input_regs_2_a6; // @[RegsRouter.scala 25:33:@40.6]
  assign _T_1002 = io_input_regs_1_a7 | io_input_regs_2_a7; // @[RegsRouter.scala 26:33:@42.6]
  assign _T_1003 = io_input_regs_1_s2 | io_input_regs_2_s2; // @[RegsRouter.scala 27:33:@44.6]
  assign _T_1004 = io_input_regs_1_s3 | io_input_regs_2_s3; // @[RegsRouter.scala 28:33:@46.6]
  assign _T_1005 = io_input_regs_1_s4 | io_input_regs_2_s4; // @[RegsRouter.scala 29:33:@48.6]
  assign _T_1006 = io_input_regs_1_s5 | io_input_regs_2_s5; // @[RegsRouter.scala 30:33:@50.6]
  assign _T_1007 = io_input_regs_1_s6 | io_input_regs_2_s6; // @[RegsRouter.scala 31:33:@52.6]
  assign _T_1008 = io_input_regs_1_s7 | io_input_regs_2_s7; // @[RegsRouter.scala 32:33:@54.6]
  assign _T_1009 = io_input_regs_1_s8 | io_input_regs_2_s8; // @[RegsRouter.scala 33:33:@56.6]
  assign _T_1010 = io_input_regs_1_s9 | io_input_regs_2_s9; // @[RegsRouter.scala 34:33:@58.6]
  assign _T_1011 = io_input_regs_1_s10 | io_input_regs_2_s10; // @[RegsRouter.scala 35:35:@60.6]
  assign _T_1012 = io_input_regs_1_s11 | io_input_regs_2_s11; // @[RegsRouter.scala 36:35:@62.6]
  assign _T_1013 = io_input_regs_1_t3 | io_input_regs_2_t3; // @[RegsRouter.scala 37:33:@64.6]
  assign _T_1014 = io_input_regs_1_t4 | io_input_regs_2_t4; // @[RegsRouter.scala 38:33:@66.6]
  assign _T_1015 = io_input_regs_1_t5 | io_input_regs_2_t5; // @[RegsRouter.scala 39:33:@68.6]
  assign _T_1016 = io_input_regs_1_t6 | io_input_regs_2_t6; // @[RegsRouter.scala 40:33:@70.6]
  assign _T_1017 = io_input_regs_1_pc | io_input_regs_2_pc; // @[RegsRouter.scala 41:33:@72.6]
  assign _T_1018 = io_input_regs_1_interrupt | io_input_regs_2_interrupt; // @[RegsRouter.scala 42:47:@74.6]
  assign _T_1019 = io_input_regs_1_interrupt_cause | io_input_regs_2_interrupt_cause; // @[RegsRouter.scala 43:59:@76.6]
  assign _T_1020 = io_input_regs_1_time | io_input_regs_2_time; // @[RegsRouter.scala 44:37:@78.6]
  assign _T_1021 = io_input_regs_1_debug | io_input_regs_2_debug; // @[RegsRouter.scala 45:39:@80.6]
  assign _T_1022 = io_input_regs_1_isa | io_input_regs_2_isa; // @[RegsRouter.scala 46:35:@82.6]
  assign _T_1023 = io_input_regs_1_sd | io_input_regs_2_sd; // @[RegsRouter.scala 47:33:@84.6]
  assign _T_1024 = io_input_regs_1_sd_rv32 | io_input_regs_2_sd_rv32; // @[RegsRouter.scala 48:43:@86.6]
  assign _T_1025 = io_input_regs_1_mpp | io_input_regs_2_mpp; // @[RegsRouter.scala 49:35:@88.6]
  assign _T_1026 = io_input_regs_1_spp | io_input_regs_2_spp; // @[RegsRouter.scala 50:35:@90.6]
  assign _T_1027 = io_input_regs_1_mpie | io_input_regs_2_mpie; // @[RegsRouter.scala 51:37:@92.6]
  assign _T_1028 = io_input_regs_1_mie | io_input_regs_2_mie; // @[RegsRouter.scala 52:35:@94.6]
  assign _T_1029 = io_input_regs_1_evec | io_input_regs_2_evec; // @[RegsRouter.scala 53:37:@96.6]
  assign _T_1030 = io_input_regs_1_ra | io_input_regs_1_ra; // @[RegsRouter.scala 10:33:@98.6]
  assign _T_1031 = io_input_regs_1_sp | io_input_regs_1_sp; // @[RegsRouter.scala 11:33:@100.6]
  assign _T_1032 = io_input_regs_1_gp | io_input_regs_1_gp; // @[RegsRouter.scala 12:33:@102.6]
  assign _T_1033 = io_input_regs_1_tp | io_input_regs_1_tp; // @[RegsRouter.scala 13:33:@104.6]
  assign _T_1034 = io_input_regs_1_t0 | io_input_regs_1_t0; // @[RegsRouter.scala 14:33:@106.6]
  assign _T_1035 = io_input_regs_1_t1 | io_input_regs_1_t1; // @[RegsRouter.scala 15:33:@108.6]
  assign _T_1036 = io_input_regs_1_t2 | io_input_regs_1_t2; // @[RegsRouter.scala 16:33:@110.6]
  assign _T_1037 = io_input_regs_1_fp | io_input_regs_1_fp; // @[RegsRouter.scala 17:33:@112.6]
  assign _T_1038 = io_input_regs_1_s1 | io_input_regs_1_s1; // @[RegsRouter.scala 18:33:@114.6]
  assign _T_1039 = io_input_regs_1_a0 | io_input_regs_1_a0; // @[RegsRouter.scala 19:33:@116.6]
  assign _T_1040 = io_input_regs_1_a1 | io_input_regs_1_a1; // @[RegsRouter.scala 20:33:@118.6]
  assign _T_1041 = io_input_regs_1_a2 | io_input_regs_1_a2; // @[RegsRouter.scala 21:33:@120.6]
  assign _T_1042 = io_input_regs_1_a3 | io_input_regs_1_a3; // @[RegsRouter.scala 22:33:@122.6]
  assign _T_1043 = io_input_regs_1_a4 | io_input_regs_1_a4; // @[RegsRouter.scala 23:33:@124.6]
  assign _T_1044 = io_input_regs_1_a5 | io_input_regs_1_a5; // @[RegsRouter.scala 24:33:@126.6]
  assign _T_1045 = io_input_regs_1_a6 | io_input_regs_1_a6; // @[RegsRouter.scala 25:33:@128.6]
  assign _T_1046 = io_input_regs_1_a7 | io_input_regs_1_a7; // @[RegsRouter.scala 26:33:@130.6]
  assign _T_1047 = io_input_regs_1_s2 | io_input_regs_1_s2; // @[RegsRouter.scala 27:33:@132.6]
  assign _T_1048 = io_input_regs_1_s3 | io_input_regs_1_s3; // @[RegsRouter.scala 28:33:@134.6]
  assign _T_1049 = io_input_regs_1_s4 | io_input_regs_1_s4; // @[RegsRouter.scala 29:33:@136.6]
  assign _T_1050 = io_input_regs_1_s5 | io_input_regs_1_s5; // @[RegsRouter.scala 30:33:@138.6]
  assign _T_1051 = io_input_regs_1_s6 | io_input_regs_1_s6; // @[RegsRouter.scala 31:33:@140.6]
  assign _T_1052 = io_input_regs_1_s7 | io_input_regs_1_s7; // @[RegsRouter.scala 32:33:@142.6]
  assign _T_1053 = io_input_regs_1_s8 | io_input_regs_1_s8; // @[RegsRouter.scala 33:33:@144.6]
  assign _T_1054 = io_input_regs_1_s9 | io_input_regs_1_s9; // @[RegsRouter.scala 34:33:@146.6]
  assign _T_1055 = io_input_regs_1_s10 | io_input_regs_1_s10; // @[RegsRouter.scala 35:35:@148.6]
  assign _T_1056 = io_input_regs_1_s11 | io_input_regs_1_s11; // @[RegsRouter.scala 36:35:@150.6]
  assign _T_1057 = io_input_regs_1_t3 | io_input_regs_1_t3; // @[RegsRouter.scala 37:33:@152.6]
  assign _T_1058 = io_input_regs_1_t4 | io_input_regs_1_t4; // @[RegsRouter.scala 38:33:@154.6]
  assign _T_1059 = io_input_regs_1_t5 | io_input_regs_1_t5; // @[RegsRouter.scala 39:33:@156.6]
  assign _T_1060 = io_input_regs_1_t6 | io_input_regs_1_t6; // @[RegsRouter.scala 40:33:@158.6]
  assign _T_1061 = io_input_regs_1_pc | io_input_regs_1_pc; // @[RegsRouter.scala 41:33:@160.6]
  assign _T_1062 = io_input_regs_1_interrupt | io_input_regs_1_interrupt; // @[RegsRouter.scala 42:47:@162.6]
  assign _T_1063 = io_input_regs_1_interrupt_cause | io_input_regs_1_interrupt_cause; // @[RegsRouter.scala 43:59:@164.6]
  assign _T_1064 = io_input_regs_1_time | io_input_regs_1_time; // @[RegsRouter.scala 44:37:@166.6]
  assign _T_1065 = io_input_regs_1_debug | io_input_regs_1_debug; // @[RegsRouter.scala 45:39:@168.6]
  assign _T_1066 = io_input_regs_1_isa | io_input_regs_1_isa; // @[RegsRouter.scala 46:35:@170.6]
  assign _T_1067 = io_input_regs_1_sd | io_input_regs_1_sd; // @[RegsRouter.scala 47:33:@172.6]
  assign _T_1068 = io_input_regs_1_sd_rv32 | io_input_regs_1_sd_rv32; // @[RegsRouter.scala 48:43:@174.6]
  assign _T_1069 = io_input_regs_1_mpp | io_input_regs_1_mpp; // @[RegsRouter.scala 49:35:@176.6]
  assign _T_1070 = io_input_regs_1_spp | io_input_regs_1_spp; // @[RegsRouter.scala 50:35:@178.6]
  assign _T_1071 = io_input_regs_1_mpie | io_input_regs_1_mpie; // @[RegsRouter.scala 51:37:@180.6]
  assign _T_1072 = io_input_regs_1_mie | io_input_regs_1_mie; // @[RegsRouter.scala 52:35:@182.6]
  assign _T_1073 = io_input_regs_1_evec | io_input_regs_1_evec; // @[RegsRouter.scala 53:37:@184.6]
  assign _T_1074 = io_input_regs_2_ra | io_input_regs_2_ra; // @[RegsRouter.scala 10:33:@186.6]
  assign _T_1075 = io_input_regs_2_sp | io_input_regs_2_sp; // @[RegsRouter.scala 11:33:@188.6]
  assign _T_1076 = io_input_regs_2_gp | io_input_regs_2_gp; // @[RegsRouter.scala 12:33:@190.6]
  assign _T_1077 = io_input_regs_2_tp | io_input_regs_2_tp; // @[RegsRouter.scala 13:33:@192.6]
  assign _T_1078 = io_input_regs_2_t0 | io_input_regs_2_t0; // @[RegsRouter.scala 14:33:@194.6]
  assign _T_1079 = io_input_regs_2_t1 | io_input_regs_2_t1; // @[RegsRouter.scala 15:33:@196.6]
  assign _T_1080 = io_input_regs_2_t2 | io_input_regs_2_t2; // @[RegsRouter.scala 16:33:@198.6]
  assign _T_1081 = io_input_regs_2_fp | io_input_regs_2_fp; // @[RegsRouter.scala 17:33:@200.6]
  assign _T_1082 = io_input_regs_2_s1 | io_input_regs_2_s1; // @[RegsRouter.scala 18:33:@202.6]
  assign _T_1083 = io_input_regs_2_a0 | io_input_regs_2_a0; // @[RegsRouter.scala 19:33:@204.6]
  assign _T_1084 = io_input_regs_2_a1 | io_input_regs_2_a1; // @[RegsRouter.scala 20:33:@206.6]
  assign _T_1085 = io_input_regs_2_a2 | io_input_regs_2_a2; // @[RegsRouter.scala 21:33:@208.6]
  assign _T_1086 = io_input_regs_2_a3 | io_input_regs_2_a3; // @[RegsRouter.scala 22:33:@210.6]
  assign _T_1087 = io_input_regs_2_a4 | io_input_regs_2_a4; // @[RegsRouter.scala 23:33:@212.6]
  assign _T_1088 = io_input_regs_2_a5 | io_input_regs_2_a5; // @[RegsRouter.scala 24:33:@214.6]
  assign _T_1089 = io_input_regs_2_a6 | io_input_regs_2_a6; // @[RegsRouter.scala 25:33:@216.6]
  assign _T_1090 = io_input_regs_2_a7 | io_input_regs_2_a7; // @[RegsRouter.scala 26:33:@218.6]
  assign _T_1091 = io_input_regs_2_s2 | io_input_regs_2_s2; // @[RegsRouter.scala 27:33:@220.6]
  assign _T_1092 = io_input_regs_2_s3 | io_input_regs_2_s3; // @[RegsRouter.scala 28:33:@222.6]
  assign _T_1093 = io_input_regs_2_s4 | io_input_regs_2_s4; // @[RegsRouter.scala 29:33:@224.6]
  assign _T_1094 = io_input_regs_2_s5 | io_input_regs_2_s5; // @[RegsRouter.scala 30:33:@226.6]
  assign _T_1095 = io_input_regs_2_s6 | io_input_regs_2_s6; // @[RegsRouter.scala 31:33:@228.6]
  assign _T_1096 = io_input_regs_2_s7 | io_input_regs_2_s7; // @[RegsRouter.scala 32:33:@230.6]
  assign _T_1097 = io_input_regs_2_s8 | io_input_regs_2_s8; // @[RegsRouter.scala 33:33:@232.6]
  assign _T_1098 = io_input_regs_2_s9 | io_input_regs_2_s9; // @[RegsRouter.scala 34:33:@234.6]
  assign _T_1099 = io_input_regs_2_s10 | io_input_regs_2_s10; // @[RegsRouter.scala 35:35:@236.6]
  assign _T_1100 = io_input_regs_2_s11 | io_input_regs_2_s11; // @[RegsRouter.scala 36:35:@238.6]
  assign _T_1101 = io_input_regs_2_t3 | io_input_regs_2_t3; // @[RegsRouter.scala 37:33:@240.6]
  assign _T_1102 = io_input_regs_2_t4 | io_input_regs_2_t4; // @[RegsRouter.scala 38:33:@242.6]
  assign _T_1103 = io_input_regs_2_t5 | io_input_regs_2_t5; // @[RegsRouter.scala 39:33:@244.6]
  assign _T_1104 = io_input_regs_2_t6 | io_input_regs_2_t6; // @[RegsRouter.scala 40:33:@246.6]
  assign _T_1105 = io_input_regs_2_pc | io_input_regs_2_pc; // @[RegsRouter.scala 41:33:@248.6]
  assign _T_1106 = io_input_regs_2_interrupt | io_input_regs_2_interrupt; // @[RegsRouter.scala 42:47:@250.6]
  assign _T_1107 = io_input_regs_2_interrupt_cause | io_input_regs_2_interrupt_cause; // @[RegsRouter.scala 43:59:@252.6]
  assign _T_1108 = io_input_regs_2_time | io_input_regs_2_time; // @[RegsRouter.scala 44:37:@254.6]
  assign _T_1109 = io_input_regs_2_debug | io_input_regs_2_debug; // @[RegsRouter.scala 45:39:@256.6]
  assign _T_1110 = io_input_regs_2_isa | io_input_regs_2_isa; // @[RegsRouter.scala 46:35:@258.6]
  assign _T_1111 = io_input_regs_2_sd | io_input_regs_2_sd; // @[RegsRouter.scala 47:33:@260.6]
  assign _T_1112 = io_input_regs_2_sd_rv32 | io_input_regs_2_sd_rv32; // @[RegsRouter.scala 48:43:@262.6]
  assign _T_1113 = io_input_regs_2_mpp | io_input_regs_2_mpp; // @[RegsRouter.scala 49:35:@264.6]
  assign _T_1114 = io_input_regs_2_spp | io_input_regs_2_spp; // @[RegsRouter.scala 50:35:@266.6]
  assign _T_1115 = io_input_regs_2_mpie | io_input_regs_2_mpie; // @[RegsRouter.scala 51:37:@268.6]
  assign _T_1116 = io_input_regs_2_mie | io_input_regs_2_mie; // @[RegsRouter.scala 52:35:@270.6]
  assign _T_1117 = io_input_regs_2_evec | io_input_regs_2_evec; // @[RegsRouter.scala 53:37:@272.6]
  assign _T_1118 = io_selector == 3'h2; // @[RegsRouter.scala 73:26:@276.6]
  assign _T_1119 = io_input_regs_0_ra | io_input_regs_0_ra; // @[RegsRouter.scala 10:33:@278.8]
  assign _T_1120 = io_input_regs_0_sp | io_input_regs_0_sp; // @[RegsRouter.scala 11:33:@280.8]
  assign _T_1121 = io_input_regs_0_gp | io_input_regs_0_gp; // @[RegsRouter.scala 12:33:@282.8]
  assign _T_1122 = io_input_regs_0_tp | io_input_regs_0_tp; // @[RegsRouter.scala 13:33:@284.8]
  assign _T_1123 = io_input_regs_0_t0 | io_input_regs_0_t0; // @[RegsRouter.scala 14:33:@286.8]
  assign _T_1124 = io_input_regs_0_t1 | io_input_regs_0_t1; // @[RegsRouter.scala 15:33:@288.8]
  assign _T_1125 = io_input_regs_0_t2 | io_input_regs_0_t2; // @[RegsRouter.scala 16:33:@290.8]
  assign _T_1126 = io_input_regs_0_fp | io_input_regs_0_fp; // @[RegsRouter.scala 17:33:@292.8]
  assign _T_1127 = io_input_regs_0_s1 | io_input_regs_0_s1; // @[RegsRouter.scala 18:33:@294.8]
  assign _T_1128 = io_input_regs_0_a0 | io_input_regs_0_a0; // @[RegsRouter.scala 19:33:@296.8]
  assign _T_1129 = io_input_regs_0_a1 | io_input_regs_0_a1; // @[RegsRouter.scala 20:33:@298.8]
  assign _T_1130 = io_input_regs_0_a2 | io_input_regs_0_a2; // @[RegsRouter.scala 21:33:@300.8]
  assign _T_1131 = io_input_regs_0_a3 | io_input_regs_0_a3; // @[RegsRouter.scala 22:33:@302.8]
  assign _T_1132 = io_input_regs_0_a4 | io_input_regs_0_a4; // @[RegsRouter.scala 23:33:@304.8]
  assign _T_1133 = io_input_regs_0_a5 | io_input_regs_0_a5; // @[RegsRouter.scala 24:33:@306.8]
  assign _T_1134 = io_input_regs_0_a6 | io_input_regs_0_a6; // @[RegsRouter.scala 25:33:@308.8]
  assign _T_1135 = io_input_regs_0_a7 | io_input_regs_0_a7; // @[RegsRouter.scala 26:33:@310.8]
  assign _T_1136 = io_input_regs_0_s2 | io_input_regs_0_s2; // @[RegsRouter.scala 27:33:@312.8]
  assign _T_1137 = io_input_regs_0_s3 | io_input_regs_0_s3; // @[RegsRouter.scala 28:33:@314.8]
  assign _T_1138 = io_input_regs_0_s4 | io_input_regs_0_s4; // @[RegsRouter.scala 29:33:@316.8]
  assign _T_1139 = io_input_regs_0_s5 | io_input_regs_0_s5; // @[RegsRouter.scala 30:33:@318.8]
  assign _T_1140 = io_input_regs_0_s6 | io_input_regs_0_s6; // @[RegsRouter.scala 31:33:@320.8]
  assign _T_1141 = io_input_regs_0_s7 | io_input_regs_0_s7; // @[RegsRouter.scala 32:33:@322.8]
  assign _T_1142 = io_input_regs_0_s8 | io_input_regs_0_s8; // @[RegsRouter.scala 33:33:@324.8]
  assign _T_1143 = io_input_regs_0_s9 | io_input_regs_0_s9; // @[RegsRouter.scala 34:33:@326.8]
  assign _T_1144 = io_input_regs_0_s10 | io_input_regs_0_s10; // @[RegsRouter.scala 35:35:@328.8]
  assign _T_1145 = io_input_regs_0_s11 | io_input_regs_0_s11; // @[RegsRouter.scala 36:35:@330.8]
  assign _T_1146 = io_input_regs_0_t3 | io_input_regs_0_t3; // @[RegsRouter.scala 37:33:@332.8]
  assign _T_1147 = io_input_regs_0_t4 | io_input_regs_0_t4; // @[RegsRouter.scala 38:33:@334.8]
  assign _T_1148 = io_input_regs_0_t5 | io_input_regs_0_t5; // @[RegsRouter.scala 39:33:@336.8]
  assign _T_1149 = io_input_regs_0_t6 | io_input_regs_0_t6; // @[RegsRouter.scala 40:33:@338.8]
  assign _T_1150 = io_input_regs_0_pc | io_input_regs_0_pc; // @[RegsRouter.scala 41:33:@340.8]
  assign _T_1151 = io_input_regs_0_interrupt | io_input_regs_0_interrupt; // @[RegsRouter.scala 42:47:@342.8]
  assign _T_1152 = io_input_regs_0_interrupt_cause | io_input_regs_0_interrupt_cause; // @[RegsRouter.scala 43:59:@344.8]
  assign _T_1153 = io_input_regs_0_time | io_input_regs_0_time; // @[RegsRouter.scala 44:37:@346.8]
  assign _T_1154 = io_input_regs_0_debug | io_input_regs_0_debug; // @[RegsRouter.scala 45:39:@348.8]
  assign _T_1155 = io_input_regs_0_isa | io_input_regs_0_isa; // @[RegsRouter.scala 46:35:@350.8]
  assign _T_1156 = io_input_regs_0_sd | io_input_regs_0_sd; // @[RegsRouter.scala 47:33:@352.8]
  assign _T_1157 = io_input_regs_0_sd_rv32 | io_input_regs_0_sd_rv32; // @[RegsRouter.scala 48:43:@354.8]
  assign _T_1158 = io_input_regs_0_mpp | io_input_regs_0_mpp; // @[RegsRouter.scala 49:35:@356.8]
  assign _T_1159 = io_input_regs_0_spp | io_input_regs_0_spp; // @[RegsRouter.scala 50:35:@358.8]
  assign _T_1160 = io_input_regs_0_mpie | io_input_regs_0_mpie; // @[RegsRouter.scala 51:37:@360.8]
  assign _T_1161 = io_input_regs_0_mie | io_input_regs_0_mie; // @[RegsRouter.scala 52:35:@362.8]
  assign _T_1162 = io_input_regs_0_evec | io_input_regs_0_evec; // @[RegsRouter.scala 53:37:@364.8]
  assign _T_1163 = io_input_regs_0_ra | io_input_regs_2_ra; // @[RegsRouter.scala 10:33:@366.8]
  assign _T_1164 = io_input_regs_0_sp | io_input_regs_2_sp; // @[RegsRouter.scala 11:33:@368.8]
  assign _T_1165 = io_input_regs_0_gp | io_input_regs_2_gp; // @[RegsRouter.scala 12:33:@370.8]
  assign _T_1166 = io_input_regs_0_tp | io_input_regs_2_tp; // @[RegsRouter.scala 13:33:@372.8]
  assign _T_1167 = io_input_regs_0_t0 | io_input_regs_2_t0; // @[RegsRouter.scala 14:33:@374.8]
  assign _T_1168 = io_input_regs_0_t1 | io_input_regs_2_t1; // @[RegsRouter.scala 15:33:@376.8]
  assign _T_1169 = io_input_regs_0_t2 | io_input_regs_2_t2; // @[RegsRouter.scala 16:33:@378.8]
  assign _T_1170 = io_input_regs_0_fp | io_input_regs_2_fp; // @[RegsRouter.scala 17:33:@380.8]
  assign _T_1171 = io_input_regs_0_s1 | io_input_regs_2_s1; // @[RegsRouter.scala 18:33:@382.8]
  assign _T_1172 = io_input_regs_0_a0 | io_input_regs_2_a0; // @[RegsRouter.scala 19:33:@384.8]
  assign _T_1173 = io_input_regs_0_a1 | io_input_regs_2_a1; // @[RegsRouter.scala 20:33:@386.8]
  assign _T_1174 = io_input_regs_0_a2 | io_input_regs_2_a2; // @[RegsRouter.scala 21:33:@388.8]
  assign _T_1175 = io_input_regs_0_a3 | io_input_regs_2_a3; // @[RegsRouter.scala 22:33:@390.8]
  assign _T_1176 = io_input_regs_0_a4 | io_input_regs_2_a4; // @[RegsRouter.scala 23:33:@392.8]
  assign _T_1177 = io_input_regs_0_a5 | io_input_regs_2_a5; // @[RegsRouter.scala 24:33:@394.8]
  assign _T_1178 = io_input_regs_0_a6 | io_input_regs_2_a6; // @[RegsRouter.scala 25:33:@396.8]
  assign _T_1179 = io_input_regs_0_a7 | io_input_regs_2_a7; // @[RegsRouter.scala 26:33:@398.8]
  assign _T_1180 = io_input_regs_0_s2 | io_input_regs_2_s2; // @[RegsRouter.scala 27:33:@400.8]
  assign _T_1181 = io_input_regs_0_s3 | io_input_regs_2_s3; // @[RegsRouter.scala 28:33:@402.8]
  assign _T_1182 = io_input_regs_0_s4 | io_input_regs_2_s4; // @[RegsRouter.scala 29:33:@404.8]
  assign _T_1183 = io_input_regs_0_s5 | io_input_regs_2_s5; // @[RegsRouter.scala 30:33:@406.8]
  assign _T_1184 = io_input_regs_0_s6 | io_input_regs_2_s6; // @[RegsRouter.scala 31:33:@408.8]
  assign _T_1185 = io_input_regs_0_s7 | io_input_regs_2_s7; // @[RegsRouter.scala 32:33:@410.8]
  assign _T_1186 = io_input_regs_0_s8 | io_input_regs_2_s8; // @[RegsRouter.scala 33:33:@412.8]
  assign _T_1187 = io_input_regs_0_s9 | io_input_regs_2_s9; // @[RegsRouter.scala 34:33:@414.8]
  assign _T_1188 = io_input_regs_0_s10 | io_input_regs_2_s10; // @[RegsRouter.scala 35:35:@416.8]
  assign _T_1189 = io_input_regs_0_s11 | io_input_regs_2_s11; // @[RegsRouter.scala 36:35:@418.8]
  assign _T_1190 = io_input_regs_0_t3 | io_input_regs_2_t3; // @[RegsRouter.scala 37:33:@420.8]
  assign _T_1191 = io_input_regs_0_t4 | io_input_regs_2_t4; // @[RegsRouter.scala 38:33:@422.8]
  assign _T_1192 = io_input_regs_0_t5 | io_input_regs_2_t5; // @[RegsRouter.scala 39:33:@424.8]
  assign _T_1193 = io_input_regs_0_t6 | io_input_regs_2_t6; // @[RegsRouter.scala 40:33:@426.8]
  assign _T_1194 = io_input_regs_0_pc | io_input_regs_2_pc; // @[RegsRouter.scala 41:33:@428.8]
  assign _T_1195 = io_input_regs_0_interrupt | io_input_regs_2_interrupt; // @[RegsRouter.scala 42:47:@430.8]
  assign _T_1196 = io_input_regs_0_interrupt_cause | io_input_regs_2_interrupt_cause; // @[RegsRouter.scala 43:59:@432.8]
  assign _T_1197 = io_input_regs_0_time | io_input_regs_2_time; // @[RegsRouter.scala 44:37:@434.8]
  assign _T_1198 = io_input_regs_0_debug | io_input_regs_2_debug; // @[RegsRouter.scala 45:39:@436.8]
  assign _T_1199 = io_input_regs_0_isa | io_input_regs_2_isa; // @[RegsRouter.scala 46:35:@438.8]
  assign _T_1200 = io_input_regs_0_sd | io_input_regs_2_sd; // @[RegsRouter.scala 47:33:@440.8]
  assign _T_1201 = io_input_regs_0_sd_rv32 | io_input_regs_2_sd_rv32; // @[RegsRouter.scala 48:43:@442.8]
  assign _T_1202 = io_input_regs_0_mpp | io_input_regs_2_mpp; // @[RegsRouter.scala 49:35:@444.8]
  assign _T_1203 = io_input_regs_0_spp | io_input_regs_2_spp; // @[RegsRouter.scala 50:35:@446.8]
  assign _T_1204 = io_input_regs_0_mpie | io_input_regs_2_mpie; // @[RegsRouter.scala 51:37:@448.8]
  assign _T_1205 = io_input_regs_0_mie | io_input_regs_2_mie; // @[RegsRouter.scala 52:35:@450.8]
  assign _T_1206 = io_input_regs_0_evec | io_input_regs_2_evec; // @[RegsRouter.scala 53:37:@452.8]
  assign _T_1251 = io_selector == 3'h4; // @[RegsRouter.scala 78:26:@544.8]
  assign _T_1340 = io_input_regs_0_ra | io_input_regs_1_ra; // @[RegsRouter.scala 10:33:@722.10]
  assign _T_1341 = io_input_regs_0_sp | io_input_regs_1_sp; // @[RegsRouter.scala 11:33:@724.10]
  assign _T_1342 = io_input_regs_0_gp | io_input_regs_1_gp; // @[RegsRouter.scala 12:33:@726.10]
  assign _T_1343 = io_input_regs_0_tp | io_input_regs_1_tp; // @[RegsRouter.scala 13:33:@728.10]
  assign _T_1344 = io_input_regs_0_t0 | io_input_regs_1_t0; // @[RegsRouter.scala 14:33:@730.10]
  assign _T_1345 = io_input_regs_0_t1 | io_input_regs_1_t1; // @[RegsRouter.scala 15:33:@732.10]
  assign _T_1346 = io_input_regs_0_t2 | io_input_regs_1_t2; // @[RegsRouter.scala 16:33:@734.10]
  assign _T_1347 = io_input_regs_0_fp | io_input_regs_1_fp; // @[RegsRouter.scala 17:33:@736.10]
  assign _T_1348 = io_input_regs_0_s1 | io_input_regs_1_s1; // @[RegsRouter.scala 18:33:@738.10]
  assign _T_1349 = io_input_regs_0_a0 | io_input_regs_1_a0; // @[RegsRouter.scala 19:33:@740.10]
  assign _T_1350 = io_input_regs_0_a1 | io_input_regs_1_a1; // @[RegsRouter.scala 20:33:@742.10]
  assign _T_1351 = io_input_regs_0_a2 | io_input_regs_1_a2; // @[RegsRouter.scala 21:33:@744.10]
  assign _T_1352 = io_input_regs_0_a3 | io_input_regs_1_a3; // @[RegsRouter.scala 22:33:@746.10]
  assign _T_1353 = io_input_regs_0_a4 | io_input_regs_1_a4; // @[RegsRouter.scala 23:33:@748.10]
  assign _T_1354 = io_input_regs_0_a5 | io_input_regs_1_a5; // @[RegsRouter.scala 24:33:@750.10]
  assign _T_1355 = io_input_regs_0_a6 | io_input_regs_1_a6; // @[RegsRouter.scala 25:33:@752.10]
  assign _T_1356 = io_input_regs_0_a7 | io_input_regs_1_a7; // @[RegsRouter.scala 26:33:@754.10]
  assign _T_1357 = io_input_regs_0_s2 | io_input_regs_1_s2; // @[RegsRouter.scala 27:33:@756.10]
  assign _T_1358 = io_input_regs_0_s3 | io_input_regs_1_s3; // @[RegsRouter.scala 28:33:@758.10]
  assign _T_1359 = io_input_regs_0_s4 | io_input_regs_1_s4; // @[RegsRouter.scala 29:33:@760.10]
  assign _T_1360 = io_input_regs_0_s5 | io_input_regs_1_s5; // @[RegsRouter.scala 30:33:@762.10]
  assign _T_1361 = io_input_regs_0_s6 | io_input_regs_1_s6; // @[RegsRouter.scala 31:33:@764.10]
  assign _T_1362 = io_input_regs_0_s7 | io_input_regs_1_s7; // @[RegsRouter.scala 32:33:@766.10]
  assign _T_1363 = io_input_regs_0_s8 | io_input_regs_1_s8; // @[RegsRouter.scala 33:33:@768.10]
  assign _T_1364 = io_input_regs_0_s9 | io_input_regs_1_s9; // @[RegsRouter.scala 34:33:@770.10]
  assign _T_1365 = io_input_regs_0_s10 | io_input_regs_1_s10; // @[RegsRouter.scala 35:35:@772.10]
  assign _T_1366 = io_input_regs_0_s11 | io_input_regs_1_s11; // @[RegsRouter.scala 36:35:@774.10]
  assign _T_1367 = io_input_regs_0_t3 | io_input_regs_1_t3; // @[RegsRouter.scala 37:33:@776.10]
  assign _T_1368 = io_input_regs_0_t4 | io_input_regs_1_t4; // @[RegsRouter.scala 38:33:@778.10]
  assign _T_1369 = io_input_regs_0_t5 | io_input_regs_1_t5; // @[RegsRouter.scala 39:33:@780.10]
  assign _T_1370 = io_input_regs_0_t6 | io_input_regs_1_t6; // @[RegsRouter.scala 40:33:@782.10]
  assign _T_1371 = io_input_regs_0_pc | io_input_regs_1_pc; // @[RegsRouter.scala 41:33:@784.10]
  assign _T_1372 = io_input_regs_0_interrupt | io_input_regs_1_interrupt; // @[RegsRouter.scala 42:47:@786.10]
  assign _T_1373 = io_input_regs_0_interrupt_cause | io_input_regs_1_interrupt_cause; // @[RegsRouter.scala 43:59:@788.10]
  assign _T_1374 = io_input_regs_0_time | io_input_regs_1_time; // @[RegsRouter.scala 44:37:@790.10]
  assign _T_1375 = io_input_regs_0_debug | io_input_regs_1_debug; // @[RegsRouter.scala 45:39:@792.10]
  assign _T_1376 = io_input_regs_0_isa | io_input_regs_1_isa; // @[RegsRouter.scala 46:35:@794.10]
  assign _T_1377 = io_input_regs_0_sd | io_input_regs_1_sd; // @[RegsRouter.scala 47:33:@796.10]
  assign _T_1378 = io_input_regs_0_sd_rv32 | io_input_regs_1_sd_rv32; // @[RegsRouter.scala 48:43:@798.10]
  assign _T_1379 = io_input_regs_0_mpp | io_input_regs_1_mpp; // @[RegsRouter.scala 49:35:@800.10]
  assign _T_1380 = io_input_regs_0_spp | io_input_regs_1_spp; // @[RegsRouter.scala 50:35:@802.10]
  assign _T_1381 = io_input_regs_0_mpie | io_input_regs_1_mpie; // @[RegsRouter.scala 51:37:@804.10]
  assign _T_1382 = io_input_regs_0_mie | io_input_regs_1_mie; // @[RegsRouter.scala 52:35:@806.10]
  assign _T_1383 = io_input_regs_0_evec | io_input_regs_1_evec; // @[RegsRouter.scala 53:37:@808.10]
  assign _GEN_0 = _T_1251 ? _T_1119 : _T_1119; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_1 = _T_1251 ? _T_1120 : _T_1120; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_2 = _T_1251 ? _T_1121 : _T_1121; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_3 = _T_1251 ? _T_1122 : _T_1122; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_4 = _T_1251 ? _T_1123 : _T_1123; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_5 = _T_1251 ? _T_1124 : _T_1124; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_6 = _T_1251 ? _T_1125 : _T_1125; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_7 = _T_1251 ? _T_1126 : _T_1126; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_8 = _T_1251 ? _T_1127 : _T_1127; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_9 = _T_1251 ? _T_1128 : _T_1128; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_10 = _T_1251 ? _T_1129 : _T_1129; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_11 = _T_1251 ? _T_1130 : _T_1130; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_12 = _T_1251 ? _T_1131 : _T_1131; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_13 = _T_1251 ? _T_1132 : _T_1132; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_14 = _T_1251 ? _T_1133 : _T_1133; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_15 = _T_1251 ? _T_1134 : _T_1134; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_16 = _T_1251 ? _T_1135 : _T_1135; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_17 = _T_1251 ? _T_1136 : _T_1136; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_18 = _T_1251 ? _T_1137 : _T_1137; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_19 = _T_1251 ? _T_1138 : _T_1138; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_20 = _T_1251 ? _T_1139 : _T_1139; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_21 = _T_1251 ? _T_1140 : _T_1140; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_22 = _T_1251 ? _T_1141 : _T_1141; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_23 = _T_1251 ? _T_1142 : _T_1142; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_24 = _T_1251 ? _T_1143 : _T_1143; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_25 = _T_1251 ? _T_1144 : _T_1144; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_26 = _T_1251 ? _T_1145 : _T_1145; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_27 = _T_1251 ? _T_1146 : _T_1146; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_28 = _T_1251 ? _T_1147 : _T_1147; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_29 = _T_1251 ? _T_1148 : _T_1148; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_30 = _T_1251 ? _T_1149 : _T_1149; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_31 = _T_1251 ? _T_1150 : _T_1150; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_32 = _T_1251 ? _T_1151 : _T_1151; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_33 = _T_1251 ? _T_1152 : _T_1152; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_34 = _T_1251 ? _T_1153 : _T_1153; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_35 = _T_1251 ? _T_1154 : _T_1154; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_36 = _T_1251 ? _T_1155 : _T_1155; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_37 = _T_1251 ? _T_1156 : _T_1156; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_38 = _T_1251 ? _T_1157 : _T_1157; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_39 = _T_1251 ? _T_1158 : _T_1158; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_40 = _T_1251 ? _T_1159 : _T_1159; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_41 = _T_1251 ? _T_1160 : _T_1160; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_42 = _T_1251 ? _T_1161 : _T_1161; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_43 = _T_1251 ? _T_1162 : _T_1162; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_44 = _T_1251 ? _T_1030 : _T_1030; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_45 = _T_1251 ? _T_1031 : _T_1031; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_46 = _T_1251 ? _T_1032 : _T_1032; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_47 = _T_1251 ? _T_1033 : _T_1033; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_48 = _T_1251 ? _T_1034 : _T_1034; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_49 = _T_1251 ? _T_1035 : _T_1035; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_50 = _T_1251 ? _T_1036 : _T_1036; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_51 = _T_1251 ? _T_1037 : _T_1037; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_52 = _T_1251 ? _T_1038 : _T_1038; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_53 = _T_1251 ? _T_1039 : _T_1039; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_54 = _T_1251 ? _T_1040 : _T_1040; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_55 = _T_1251 ? _T_1041 : _T_1041; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_56 = _T_1251 ? _T_1042 : _T_1042; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_57 = _T_1251 ? _T_1043 : _T_1043; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_58 = _T_1251 ? _T_1044 : _T_1044; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_59 = _T_1251 ? _T_1045 : _T_1045; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_60 = _T_1251 ? _T_1046 : _T_1046; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_61 = _T_1251 ? _T_1047 : _T_1047; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_62 = _T_1251 ? _T_1048 : _T_1048; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_63 = _T_1251 ? _T_1049 : _T_1049; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_64 = _T_1251 ? _T_1050 : _T_1050; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_65 = _T_1251 ? _T_1051 : _T_1051; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_66 = _T_1251 ? _T_1052 : _T_1052; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_67 = _T_1251 ? _T_1053 : _T_1053; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_68 = _T_1251 ? _T_1054 : _T_1054; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_69 = _T_1251 ? _T_1055 : _T_1055; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_70 = _T_1251 ? _T_1056 : _T_1056; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_71 = _T_1251 ? _T_1057 : _T_1057; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_72 = _T_1251 ? _T_1058 : _T_1058; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_73 = _T_1251 ? _T_1059 : _T_1059; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_74 = _T_1251 ? _T_1060 : _T_1060; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_75 = _T_1251 ? _T_1061 : _T_1061; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_76 = _T_1251 ? _T_1062 : _T_1062; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_77 = _T_1251 ? _T_1063 : _T_1063; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_78 = _T_1251 ? _T_1064 : _T_1064; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_79 = _T_1251 ? _T_1065 : _T_1065; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_80 = _T_1251 ? _T_1066 : _T_1066; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_81 = _T_1251 ? _T_1067 : _T_1067; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_82 = _T_1251 ? _T_1068 : _T_1068; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_83 = _T_1251 ? _T_1069 : _T_1069; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_84 = _T_1251 ? _T_1070 : _T_1070; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_85 = _T_1251 ? _T_1071 : _T_1071; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_86 = _T_1251 ? _T_1072 : _T_1072; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_87 = _T_1251 ? _T_1073 : _T_1073; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_88 = _T_1251 ? _T_1340 : _T_1074; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_89 = _T_1251 ? _T_1341 : _T_1075; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_90 = _T_1251 ? _T_1342 : _T_1076; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_91 = _T_1251 ? _T_1343 : _T_1077; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_92 = _T_1251 ? _T_1344 : _T_1078; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_93 = _T_1251 ? _T_1345 : _T_1079; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_94 = _T_1251 ? _T_1346 : _T_1080; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_95 = _T_1251 ? _T_1347 : _T_1081; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_96 = _T_1251 ? _T_1348 : _T_1082; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_97 = _T_1251 ? _T_1349 : _T_1083; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_98 = _T_1251 ? _T_1350 : _T_1084; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_99 = _T_1251 ? _T_1351 : _T_1085; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_100 = _T_1251 ? _T_1352 : _T_1086; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_101 = _T_1251 ? _T_1353 : _T_1087; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_102 = _T_1251 ? _T_1354 : _T_1088; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_103 = _T_1251 ? _T_1355 : _T_1089; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_104 = _T_1251 ? _T_1356 : _T_1090; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_105 = _T_1251 ? _T_1357 : _T_1091; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_106 = _T_1251 ? _T_1358 : _T_1092; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_107 = _T_1251 ? _T_1359 : _T_1093; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_108 = _T_1251 ? _T_1360 : _T_1094; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_109 = _T_1251 ? _T_1361 : _T_1095; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_110 = _T_1251 ? _T_1362 : _T_1096; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_111 = _T_1251 ? _T_1363 : _T_1097; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_112 = _T_1251 ? _T_1364 : _T_1098; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_113 = _T_1251 ? _T_1365 : _T_1099; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_114 = _T_1251 ? _T_1366 : _T_1100; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_115 = _T_1251 ? _T_1367 : _T_1101; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_116 = _T_1251 ? _T_1368 : _T_1102; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_117 = _T_1251 ? _T_1369 : _T_1103; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_118 = _T_1251 ? _T_1370 : _T_1104; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_119 = _T_1251 ? _T_1371 : _T_1105; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_120 = _T_1251 ? _T_1372 : _T_1106; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_121 = _T_1251 ? _T_1373 : _T_1107; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_122 = _T_1251 ? _T_1374 : _T_1108; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_123 = _T_1251 ? _T_1375 : _T_1109; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_124 = _T_1251 ? _T_1376 : _T_1110; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_125 = _T_1251 ? _T_1377 : _T_1111; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_126 = _T_1251 ? _T_1378 : _T_1112; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_127 = _T_1251 ? _T_1379 : _T_1113; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_128 = _T_1251 ? _T_1380 : _T_1114; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_129 = _T_1251 ? _T_1381 : _T_1115; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_130 = _T_1251 ? _T_1382 : _T_1116; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_131 = _T_1251 ? _T_1383 : _T_1117; // @[RegsRouter.scala 78:44:@545.8]
  assign _GEN_132 = _T_1118 ? _T_1119 : _GEN_0; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_133 = _T_1118 ? _T_1120 : _GEN_1; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_134 = _T_1118 ? _T_1121 : _GEN_2; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_135 = _T_1118 ? _T_1122 : _GEN_3; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_136 = _T_1118 ? _T_1123 : _GEN_4; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_137 = _T_1118 ? _T_1124 : _GEN_5; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_138 = _T_1118 ? _T_1125 : _GEN_6; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_139 = _T_1118 ? _T_1126 : _GEN_7; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_140 = _T_1118 ? _T_1127 : _GEN_8; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_141 = _T_1118 ? _T_1128 : _GEN_9; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_142 = _T_1118 ? _T_1129 : _GEN_10; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_143 = _T_1118 ? _T_1130 : _GEN_11; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_144 = _T_1118 ? _T_1131 : _GEN_12; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_145 = _T_1118 ? _T_1132 : _GEN_13; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_146 = _T_1118 ? _T_1133 : _GEN_14; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_147 = _T_1118 ? _T_1134 : _GEN_15; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_148 = _T_1118 ? _T_1135 : _GEN_16; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_149 = _T_1118 ? _T_1136 : _GEN_17; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_150 = _T_1118 ? _T_1137 : _GEN_18; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_151 = _T_1118 ? _T_1138 : _GEN_19; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_152 = _T_1118 ? _T_1139 : _GEN_20; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_153 = _T_1118 ? _T_1140 : _GEN_21; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_154 = _T_1118 ? _T_1141 : _GEN_22; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_155 = _T_1118 ? _T_1142 : _GEN_23; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_156 = _T_1118 ? _T_1143 : _GEN_24; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_157 = _T_1118 ? _T_1144 : _GEN_25; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_158 = _T_1118 ? _T_1145 : _GEN_26; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_159 = _T_1118 ? _T_1146 : _GEN_27; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_160 = _T_1118 ? _T_1147 : _GEN_28; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_161 = _T_1118 ? _T_1148 : _GEN_29; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_162 = _T_1118 ? _T_1149 : _GEN_30; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_163 = _T_1118 ? _T_1150 : _GEN_31; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_164 = _T_1118 ? _T_1151 : _GEN_32; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_165 = _T_1118 ? _T_1152 : _GEN_33; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_166 = _T_1118 ? _T_1153 : _GEN_34; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_167 = _T_1118 ? _T_1154 : _GEN_35; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_168 = _T_1118 ? _T_1155 : _GEN_36; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_169 = _T_1118 ? _T_1156 : _GEN_37; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_170 = _T_1118 ? _T_1157 : _GEN_38; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_171 = _T_1118 ? _T_1158 : _GEN_39; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_172 = _T_1118 ? _T_1159 : _GEN_40; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_173 = _T_1118 ? _T_1160 : _GEN_41; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_174 = _T_1118 ? _T_1161 : _GEN_42; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_175 = _T_1118 ? _T_1162 : _GEN_43; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_176 = _T_1118 ? _T_1163 : _GEN_44; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_177 = _T_1118 ? _T_1164 : _GEN_45; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_178 = _T_1118 ? _T_1165 : _GEN_46; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_179 = _T_1118 ? _T_1166 : _GEN_47; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_180 = _T_1118 ? _T_1167 : _GEN_48; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_181 = _T_1118 ? _T_1168 : _GEN_49; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_182 = _T_1118 ? _T_1169 : _GEN_50; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_183 = _T_1118 ? _T_1170 : _GEN_51; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_184 = _T_1118 ? _T_1171 : _GEN_52; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_185 = _T_1118 ? _T_1172 : _GEN_53; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_186 = _T_1118 ? _T_1173 : _GEN_54; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_187 = _T_1118 ? _T_1174 : _GEN_55; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_188 = _T_1118 ? _T_1175 : _GEN_56; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_189 = _T_1118 ? _T_1176 : _GEN_57; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_190 = _T_1118 ? _T_1177 : _GEN_58; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_191 = _T_1118 ? _T_1178 : _GEN_59; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_192 = _T_1118 ? _T_1179 : _GEN_60; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_193 = _T_1118 ? _T_1180 : _GEN_61; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_194 = _T_1118 ? _T_1181 : _GEN_62; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_195 = _T_1118 ? _T_1182 : _GEN_63; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_196 = _T_1118 ? _T_1183 : _GEN_64; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_197 = _T_1118 ? _T_1184 : _GEN_65; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_198 = _T_1118 ? _T_1185 : _GEN_66; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_199 = _T_1118 ? _T_1186 : _GEN_67; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_200 = _T_1118 ? _T_1187 : _GEN_68; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_201 = _T_1118 ? _T_1188 : _GEN_69; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_202 = _T_1118 ? _T_1189 : _GEN_70; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_203 = _T_1118 ? _T_1190 : _GEN_71; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_204 = _T_1118 ? _T_1191 : _GEN_72; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_205 = _T_1118 ? _T_1192 : _GEN_73; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_206 = _T_1118 ? _T_1193 : _GEN_74; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_207 = _T_1118 ? _T_1194 : _GEN_75; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_208 = _T_1118 ? _T_1195 : _GEN_76; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_209 = _T_1118 ? _T_1196 : _GEN_77; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_210 = _T_1118 ? _T_1197 : _GEN_78; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_211 = _T_1118 ? _T_1198 : _GEN_79; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_212 = _T_1118 ? _T_1199 : _GEN_80; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_213 = _T_1118 ? _T_1200 : _GEN_81; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_214 = _T_1118 ? _T_1201 : _GEN_82; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_215 = _T_1118 ? _T_1202 : _GEN_83; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_216 = _T_1118 ? _T_1203 : _GEN_84; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_217 = _T_1118 ? _T_1204 : _GEN_85; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_218 = _T_1118 ? _T_1205 : _GEN_86; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_219 = _T_1118 ? _T_1206 : _GEN_87; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_220 = _T_1118 ? _T_1074 : _GEN_88; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_221 = _T_1118 ? _T_1075 : _GEN_89; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_222 = _T_1118 ? _T_1076 : _GEN_90; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_223 = _T_1118 ? _T_1077 : _GEN_91; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_224 = _T_1118 ? _T_1078 : _GEN_92; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_225 = _T_1118 ? _T_1079 : _GEN_93; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_226 = _T_1118 ? _T_1080 : _GEN_94; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_227 = _T_1118 ? _T_1081 : _GEN_95; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_228 = _T_1118 ? _T_1082 : _GEN_96; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_229 = _T_1118 ? _T_1083 : _GEN_97; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_230 = _T_1118 ? _T_1084 : _GEN_98; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_231 = _T_1118 ? _T_1085 : _GEN_99; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_232 = _T_1118 ? _T_1086 : _GEN_100; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_233 = _T_1118 ? _T_1087 : _GEN_101; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_234 = _T_1118 ? _T_1088 : _GEN_102; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_235 = _T_1118 ? _T_1089 : _GEN_103; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_236 = _T_1118 ? _T_1090 : _GEN_104; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_237 = _T_1118 ? _T_1091 : _GEN_105; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_238 = _T_1118 ? _T_1092 : _GEN_106; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_239 = _T_1118 ? _T_1093 : _GEN_107; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_240 = _T_1118 ? _T_1094 : _GEN_108; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_241 = _T_1118 ? _T_1095 : _GEN_109; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_242 = _T_1118 ? _T_1096 : _GEN_110; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_243 = _T_1118 ? _T_1097 : _GEN_111; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_244 = _T_1118 ? _T_1098 : _GEN_112; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_245 = _T_1118 ? _T_1099 : _GEN_113; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_246 = _T_1118 ? _T_1100 : _GEN_114; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_247 = _T_1118 ? _T_1101 : _GEN_115; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_248 = _T_1118 ? _T_1102 : _GEN_116; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_249 = _T_1118 ? _T_1103 : _GEN_117; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_250 = _T_1118 ? _T_1104 : _GEN_118; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_251 = _T_1118 ? _T_1105 : _GEN_119; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_252 = _T_1118 ? _T_1106 : _GEN_120; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_253 = _T_1118 ? _T_1107 : _GEN_121; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_254 = _T_1118 ? _T_1108 : _GEN_122; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_255 = _T_1118 ? _T_1109 : _GEN_123; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_256 = _T_1118 ? _T_1110 : _GEN_124; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_257 = _T_1118 ? _T_1111 : _GEN_125; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_258 = _T_1118 ? _T_1112 : _GEN_126; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_259 = _T_1118 ? _T_1113 : _GEN_127; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_260 = _T_1118 ? _T_1114 : _GEN_128; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_261 = _T_1118 ? _T_1115 : _GEN_129; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_262 = _T_1118 ? _T_1116 : _GEN_130; // @[RegsRouter.scala 73:44:@277.6]
  assign _GEN_263 = _T_1118 ? _T_1117 : _GEN_131; // @[RegsRouter.scala 73:44:@277.6]
  assign io_output_regs_0_ra = _T_985 ? _T_986 : _GEN_132;
  assign io_output_regs_0_sp = _T_985 ? _T_987 : _GEN_133;
  assign io_output_regs_0_gp = _T_985 ? _T_988 : _GEN_134;
  assign io_output_regs_0_tp = _T_985 ? _T_989 : _GEN_135;
  assign io_output_regs_0_t0 = _T_985 ? _T_990 : _GEN_136;
  assign io_output_regs_0_t1 = _T_985 ? _T_991 : _GEN_137;
  assign io_output_regs_0_t2 = _T_985 ? _T_992 : _GEN_138;
  assign io_output_regs_0_fp = _T_985 ? _T_993 : _GEN_139;
  assign io_output_regs_0_s1 = _T_985 ? _T_994 : _GEN_140;
  assign io_output_regs_0_a0 = _T_985 ? _T_995 : _GEN_141;
  assign io_output_regs_0_a1 = _T_985 ? _T_996 : _GEN_142;
  assign io_output_regs_0_a2 = _T_985 ? _T_997 : _GEN_143;
  assign io_output_regs_0_a3 = _T_985 ? _T_998 : _GEN_144;
  assign io_output_regs_0_a4 = _T_985 ? _T_999 : _GEN_145;
  assign io_output_regs_0_a5 = _T_985 ? _T_1000 : _GEN_146;
  assign io_output_regs_0_a6 = _T_985 ? _T_1001 : _GEN_147;
  assign io_output_regs_0_a7 = _T_985 ? _T_1002 : _GEN_148;
  assign io_output_regs_0_s2 = _T_985 ? _T_1003 : _GEN_149;
  assign io_output_regs_0_s3 = _T_985 ? _T_1004 : _GEN_150;
  assign io_output_regs_0_s4 = _T_985 ? _T_1005 : _GEN_151;
  assign io_output_regs_0_s5 = _T_985 ? _T_1006 : _GEN_152;
  assign io_output_regs_0_s6 = _T_985 ? _T_1007 : _GEN_153;
  assign io_output_regs_0_s7 = _T_985 ? _T_1008 : _GEN_154;
  assign io_output_regs_0_s8 = _T_985 ? _T_1009 : _GEN_155;
  assign io_output_regs_0_s9 = _T_985 ? _T_1010 : _GEN_156;
  assign io_output_regs_0_s10 = _T_985 ? _T_1011 : _GEN_157;
  assign io_output_regs_0_s11 = _T_985 ? _T_1012 : _GEN_158;
  assign io_output_regs_0_t3 = _T_985 ? _T_1013 : _GEN_159;
  assign io_output_regs_0_t4 = _T_985 ? _T_1014 : _GEN_160;
  assign io_output_regs_0_t5 = _T_985 ? _T_1015 : _GEN_161;
  assign io_output_regs_0_t6 = _T_985 ? _T_1016 : _GEN_162;
  assign io_output_regs_0_pc = _T_985 ? _T_1017 : _GEN_163;
  assign io_output_regs_0_interrupt = _T_985 ? _T_1018 : _GEN_164;
  assign io_output_regs_0_interrupt_cause = _T_985 ? _T_1019 : _GEN_165;
  assign io_output_regs_0_time = _T_985 ? _T_1020 : _GEN_166;
  assign io_output_regs_0_debug = _T_985 ? _T_1021 : _GEN_167;
  assign io_output_regs_0_isa = _T_985 ? _T_1022 : _GEN_168;
  assign io_output_regs_0_sd = _T_985 ? _T_1023 : _GEN_169;
  assign io_output_regs_0_sd_rv32 = _T_985 ? _T_1024 : _GEN_170;
  assign io_output_regs_0_mpp = _T_985 ? _T_1025 : _GEN_171;
  assign io_output_regs_0_spp = _T_985 ? _T_1026 : _GEN_172;
  assign io_output_regs_0_mpie = _T_985 ? _T_1027 : _GEN_173;
  assign io_output_regs_0_mie = _T_985 ? _T_1028 : _GEN_174;
  assign io_output_regs_0_evec = _T_985 ? _T_1029 : _GEN_175;
  assign io_output_regs_1_ra = _T_985 ? _T_1030 : _GEN_176;
  assign io_output_regs_1_sp = _T_985 ? _T_1031 : _GEN_177;
  assign io_output_regs_1_gp = _T_985 ? _T_1032 : _GEN_178;
  assign io_output_regs_1_tp = _T_985 ? _T_1033 : _GEN_179;
  assign io_output_regs_1_t0 = _T_985 ? _T_1034 : _GEN_180;
  assign io_output_regs_1_t1 = _T_985 ? _T_1035 : _GEN_181;
  assign io_output_regs_1_t2 = _T_985 ? _T_1036 : _GEN_182;
  assign io_output_regs_1_fp = _T_985 ? _T_1037 : _GEN_183;
  assign io_output_regs_1_s1 = _T_985 ? _T_1038 : _GEN_184;
  assign io_output_regs_1_a0 = _T_985 ? _T_1039 : _GEN_185;
  assign io_output_regs_1_a1 = _T_985 ? _T_1040 : _GEN_186;
  assign io_output_regs_1_a2 = _T_985 ? _T_1041 : _GEN_187;
  assign io_output_regs_1_a3 = _T_985 ? _T_1042 : _GEN_188;
  assign io_output_regs_1_a4 = _T_985 ? _T_1043 : _GEN_189;
  assign io_output_regs_1_a5 = _T_985 ? _T_1044 : _GEN_190;
  assign io_output_regs_1_a6 = _T_985 ? _T_1045 : _GEN_191;
  assign io_output_regs_1_a7 = _T_985 ? _T_1046 : _GEN_192;
  assign io_output_regs_1_s2 = _T_985 ? _T_1047 : _GEN_193;
  assign io_output_regs_1_s3 = _T_985 ? _T_1048 : _GEN_194;
  assign io_output_regs_1_s4 = _T_985 ? _T_1049 : _GEN_195;
  assign io_output_regs_1_s5 = _T_985 ? _T_1050 : _GEN_196;
  assign io_output_regs_1_s6 = _T_985 ? _T_1051 : _GEN_197;
  assign io_output_regs_1_s7 = _T_985 ? _T_1052 : _GEN_198;
  assign io_output_regs_1_s8 = _T_985 ? _T_1053 : _GEN_199;
  assign io_output_regs_1_s9 = _T_985 ? _T_1054 : _GEN_200;
  assign io_output_regs_1_s10 = _T_985 ? _T_1055 : _GEN_201;
  assign io_output_regs_1_s11 = _T_985 ? _T_1056 : _GEN_202;
  assign io_output_regs_1_t3 = _T_985 ? _T_1057 : _GEN_203;
  assign io_output_regs_1_t4 = _T_985 ? _T_1058 : _GEN_204;
  assign io_output_regs_1_t5 = _T_985 ? _T_1059 : _GEN_205;
  assign io_output_regs_1_t6 = _T_985 ? _T_1060 : _GEN_206;
  assign io_output_regs_1_pc = _T_985 ? _T_1061 : _GEN_207;
  assign io_output_regs_1_interrupt = _T_985 ? _T_1062 : _GEN_208;
  assign io_output_regs_1_interrupt_cause = _T_985 ? _T_1063 : _GEN_209;
  assign io_output_regs_1_time = _T_985 ? _T_1064 : _GEN_210;
  assign io_output_regs_1_debug = _T_985 ? _T_1065 : _GEN_211;
  assign io_output_regs_1_isa = _T_985 ? _T_1066 : _GEN_212;
  assign io_output_regs_1_sd = _T_985 ? _T_1067 : _GEN_213;
  assign io_output_regs_1_sd_rv32 = _T_985 ? _T_1068 : _GEN_214;
  assign io_output_regs_1_mpp = _T_985 ? _T_1069 : _GEN_215;
  assign io_output_regs_1_spp = _T_985 ? _T_1070 : _GEN_216;
  assign io_output_regs_1_mpie = _T_985 ? _T_1071 : _GEN_217;
  assign io_output_regs_1_mie = _T_985 ? _T_1072 : _GEN_218;
  assign io_output_regs_1_evec = _T_985 ? _T_1073 : _GEN_219;
  assign io_output_regs_2_ra = _T_985 ? _T_1074 : _GEN_220;
  assign io_output_regs_2_sp = _T_985 ? _T_1075 : _GEN_221;
  assign io_output_regs_2_gp = _T_985 ? _T_1076 : _GEN_222;
  assign io_output_regs_2_tp = _T_985 ? _T_1077 : _GEN_223;
  assign io_output_regs_2_t0 = _T_985 ? _T_1078 : _GEN_224;
  assign io_output_regs_2_t1 = _T_985 ? _T_1079 : _GEN_225;
  assign io_output_regs_2_t2 = _T_985 ? _T_1080 : _GEN_226;
  assign io_output_regs_2_fp = _T_985 ? _T_1081 : _GEN_227;
  assign io_output_regs_2_s1 = _T_985 ? _T_1082 : _GEN_228;
  assign io_output_regs_2_a0 = _T_985 ? _T_1083 : _GEN_229;
  assign io_output_regs_2_a1 = _T_985 ? _T_1084 : _GEN_230;
  assign io_output_regs_2_a2 = _T_985 ? _T_1085 : _GEN_231;
  assign io_output_regs_2_a3 = _T_985 ? _T_1086 : _GEN_232;
  assign io_output_regs_2_a4 = _T_985 ? _T_1087 : _GEN_233;
  assign io_output_regs_2_a5 = _T_985 ? _T_1088 : _GEN_234;
  assign io_output_regs_2_a6 = _T_985 ? _T_1089 : _GEN_235;
  assign io_output_regs_2_a7 = _T_985 ? _T_1090 : _GEN_236;
  assign io_output_regs_2_s2 = _T_985 ? _T_1091 : _GEN_237;
  assign io_output_regs_2_s3 = _T_985 ? _T_1092 : _GEN_238;
  assign io_output_regs_2_s4 = _T_985 ? _T_1093 : _GEN_239;
  assign io_output_regs_2_s5 = _T_985 ? _T_1094 : _GEN_240;
  assign io_output_regs_2_s6 = _T_985 ? _T_1095 : _GEN_241;
  assign io_output_regs_2_s7 = _T_985 ? _T_1096 : _GEN_242;
  assign io_output_regs_2_s8 = _T_985 ? _T_1097 : _GEN_243;
  assign io_output_regs_2_s9 = _T_985 ? _T_1098 : _GEN_244;
  assign io_output_regs_2_s10 = _T_985 ? _T_1099 : _GEN_245;
  assign io_output_regs_2_s11 = _T_985 ? _T_1100 : _GEN_246;
  assign io_output_regs_2_t3 = _T_985 ? _T_1101 : _GEN_247;
  assign io_output_regs_2_t4 = _T_985 ? _T_1102 : _GEN_248;
  assign io_output_regs_2_t5 = _T_985 ? _T_1103 : _GEN_249;
  assign io_output_regs_2_t6 = _T_985 ? _T_1104 : _GEN_250;
  assign io_output_regs_2_pc = _T_985 ? _T_1105 : _GEN_251;
  assign io_output_regs_2_interrupt = _T_985 ? _T_1106 : _GEN_252;
  assign io_output_regs_2_interrupt_cause = _T_985 ? _T_1107 : _GEN_253;
  assign io_output_regs_2_time = _T_985 ? _T_1108 : _GEN_254;
  assign io_output_regs_2_debug = _T_985 ? _T_1109 : _GEN_255;
  assign io_output_regs_2_isa = _T_985 ? _T_1110 : _GEN_256;
  assign io_output_regs_2_sd = _T_985 ? _T_1111 : _GEN_257;
  assign io_output_regs_2_sd_rv32 = _T_985 ? _T_1112 : _GEN_258;
  assign io_output_regs_2_mpp = _T_985 ? _T_1113 : _GEN_259;
  assign io_output_regs_2_spp = _T_985 ? _T_1114 : _GEN_260;
  assign io_output_regs_2_mpie = _T_985 ? _T_1115 : _GEN_261;
  assign io_output_regs_2_mie = _T_985 ? _T_1116 : _GEN_262;
  assign io_output_regs_2_evec = _T_985 ? _T_1117 : _GEN_263;
endmodule

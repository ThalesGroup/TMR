`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module cpuRepair( // @[:@3.2]
  input   clock, // @[:@4.4]
  input   reset, // @[:@5.4]
  input   io_fault, // @[:@6.4]
  input   io_cpus_ok, // @[:@6.4]
  input   io_reset_pending, // @[:@6.4]
  output  io_ack_cpus_ok, // @[:@6.4]
  output  io_stop_cpus, // @[:@6.4]
  output  io_latch_regs, // @[:@6.4]
  output  io_reset_to_recovery, // @[:@6.4]
  output  io_reset_cpus, // @[:@6.4]
  output  io_reset_routing_logic, // @[:@6.4]
  input   io_cpu_in_interrupt // @[:@6.4]
);
  reg [2:0] state; // @[FaultDetector.scala 23:22:@8.4]
  reg [31:0] _RAND_0;
  reg  ack_cpus_ok; // @[FaultDetector.scala 25:28:@9.4]
  reg [31:0] _RAND_1;
  reg  stop_cpus; // @[FaultDetector.scala 26:26:@10.4]
  reg [31:0] _RAND_2;
  reg  latch_regs; // @[FaultDetector.scala 27:27:@11.4]
  reg [31:0] _RAND_3;
  reg  reset_to_recovery; // @[FaultDetector.scala 28:34:@12.4]
  reg [31:0] _RAND_4;
  reg  reset_cpus; // @[FaultDetector.scala 29:27:@13.4]
  reg [31:0] _RAND_5;
  reg  reset_routing_logic; // @[FaultDetector.scala 30:36:@14.4]
  reg [31:0] _RAND_6;
  wire  _T_25; // @[Conditional.scala 36:30:@15.4]
  wire [2:0] _GEN_0; // @[FaultDetector.scala 38:21:@21.6]
  wire  _T_30; // @[Conditional.scala 36:30:@26.6]
  wire  _T_33; // @[Conditional.scala 36:30:@33.8]
  wire  _T_35; // @[FaultDetector.scala 48:12:@35.10]
  wire [2:0] _GEN_1; // @[FaultDetector.scala 48:34:@36.10]
  wire  _GEN_2; // @[FaultDetector.scala 48:34:@36.10]
  wire  _T_37; // @[Conditional.scala 36:30:@42.10]
  wire  _T_39; // @[Conditional.scala 36:30:@48.12]
  wire  _T_42; // @[Conditional.scala 36:30:@55.14]
  wire [2:0] _GEN_3; // @[FaultDetector.scala 63:30:@57.16]
  wire  _T_43; // @[Conditional.scala 36:30:@62.16]
  wire  _T_45; // @[FaultDetector.scala 68:12:@64.18]
  wire [2:0] _GEN_4; // @[FaultDetector.scala 68:31:@65.18]
  wire  _GEN_5; // @[FaultDetector.scala 68:31:@65.18]
  wire  _GEN_6; // @[FaultDetector.scala 68:31:@65.18]
  wire  _T_48; // @[Conditional.scala 36:30:@72.18]
  wire  _GEN_7; // @[FaultDetector.scala 77:24:@75.20]
  wire  _GEN_8; // @[FaultDetector.scala 77:24:@75.20]
  wire [2:0] _GEN_9; // @[FaultDetector.scala 77:24:@75.20]
  wire  _GEN_10; // @[Conditional.scala 38:67:@73.18]
  wire  _GEN_11; // @[Conditional.scala 38:67:@73.18]
  wire  _GEN_12; // @[Conditional.scala 38:67:@73.18]
  wire [2:0] _GEN_13; // @[Conditional.scala 38:67:@73.18]
  wire [2:0] _GEN_14; // @[Conditional.scala 38:67:@63.16]
  wire  _GEN_15; // @[Conditional.scala 38:67:@63.16]
  wire  _GEN_16; // @[Conditional.scala 38:67:@63.16]
  wire  _GEN_17; // @[Conditional.scala 38:67:@63.16]
  wire [2:0] _GEN_18; // @[Conditional.scala 38:67:@56.14]
  wire  _GEN_19; // @[Conditional.scala 38:67:@56.14]
  wire  _GEN_20; // @[Conditional.scala 38:67:@56.14]
  wire  _GEN_21; // @[Conditional.scala 38:67:@56.14]
  wire [2:0] _GEN_22; // @[Conditional.scala 38:67:@49.12]
  wire  _GEN_23; // @[Conditional.scala 38:67:@49.12]
  wire  _GEN_24; // @[Conditional.scala 38:67:@49.12]
  wire  _GEN_25; // @[Conditional.scala 38:67:@49.12]
  wire  _GEN_26; // @[Conditional.scala 38:67:@49.12]
  wire [2:0] _GEN_27; // @[Conditional.scala 38:67:@43.10]
  wire  _GEN_28; // @[Conditional.scala 38:67:@43.10]
  wire  _GEN_29; // @[Conditional.scala 38:67:@43.10]
  wire  _GEN_30; // @[Conditional.scala 38:67:@43.10]
  wire  _GEN_31; // @[Conditional.scala 38:67:@43.10]
  wire  _GEN_32; // @[Conditional.scala 38:67:@43.10]
  wire [2:0] _GEN_33; // @[Conditional.scala 38:67:@34.8]
  wire  _GEN_34; // @[Conditional.scala 38:67:@34.8]
  wire  _GEN_35; // @[Conditional.scala 38:67:@34.8]
  wire  _GEN_36; // @[Conditional.scala 38:67:@34.8]
  wire  _GEN_37; // @[Conditional.scala 38:67:@34.8]
  wire  _GEN_38; // @[Conditional.scala 38:67:@34.8]
  wire  _GEN_39; // @[Conditional.scala 38:67:@27.6]
  wire [2:0] _GEN_40; // @[Conditional.scala 38:67:@27.6]
  wire  _GEN_41; // @[Conditional.scala 38:67:@27.6]
  wire  _GEN_42; // @[Conditional.scala 38:67:@27.6]
  wire  _GEN_43; // @[Conditional.scala 38:67:@27.6]
  wire  _GEN_44; // @[Conditional.scala 38:67:@27.6]
  wire  _GEN_45; // @[Conditional.scala 38:67:@27.6]
  wire  _GEN_46; // @[Conditional.scala 39:58:@16.4]
  wire  _GEN_47; // @[Conditional.scala 39:58:@16.4]
  wire  _GEN_48; // @[Conditional.scala 39:58:@16.4]
  wire  _GEN_49; // @[Conditional.scala 39:58:@16.4]
  wire [2:0] _GEN_50; // @[Conditional.scala 39:58:@16.4]
  wire  _GEN_51; // @[Conditional.scala 39:58:@16.4]
  wire  _GEN_52; // @[Conditional.scala 39:58:@16.4]
  assign _T_25 = 3'h0 == state; // @[Conditional.scala 36:30:@15.4]
  assign _GEN_0 = io_fault ? 3'h1 : state; // @[FaultDetector.scala 38:21:@21.6]
  assign _T_30 = 3'h1 == state; // @[Conditional.scala 36:30:@26.6]
  assign _T_33 = 3'h2 == state; // @[Conditional.scala 36:30:@33.8]
  assign _T_35 = io_cpu_in_interrupt == 1'h0; // @[FaultDetector.scala 48:12:@35.10]
  assign _GEN_1 = _T_35 ? 3'h3 : state; // @[FaultDetector.scala 48:34:@36.10]
  assign _GEN_2 = _T_35 ? 1'h1 : latch_regs; // @[FaultDetector.scala 48:34:@36.10]
  assign _T_37 = 3'h3 == state; // @[Conditional.scala 36:30:@42.10]
  assign _T_39 = 3'h4 == state; // @[Conditional.scala 36:30:@48.12]
  assign _T_42 = 3'h5 == state; // @[Conditional.scala 36:30:@55.14]
  assign _GEN_3 = io_reset_pending ? 3'h6 : state; // @[FaultDetector.scala 63:30:@57.16]
  assign _T_43 = 3'h6 == state; // @[Conditional.scala 36:30:@62.16]
  assign _T_45 = io_reset_pending == 1'h0; // @[FaultDetector.scala 68:12:@64.18]
  assign _GEN_4 = _T_45 ? 3'h7 : state; // @[FaultDetector.scala 68:31:@65.18]
  assign _GEN_5 = _T_45 ? 1'h1 : reset_routing_logic; // @[FaultDetector.scala 68:31:@65.18]
  assign _GEN_6 = _T_45 ? 1'h0 : reset_cpus; // @[FaultDetector.scala 68:31:@65.18]
  assign _T_48 = 3'h7 == state; // @[Conditional.scala 36:30:@72.18]
  assign _GEN_7 = io_cpus_ok ? 1'h0 : reset_routing_logic; // @[FaultDetector.scala 77:24:@75.20]
  assign _GEN_8 = io_cpus_ok ? 1'h1 : ack_cpus_ok; // @[FaultDetector.scala 77:24:@75.20]
  assign _GEN_9 = io_cpus_ok ? 3'h0 : state; // @[FaultDetector.scala 77:24:@75.20]
  assign _GEN_10 = _T_48 ? 1'h0 : reset_cpus; // @[Conditional.scala 38:67:@73.18]
  assign _GEN_11 = _T_48 ? _GEN_7 : reset_routing_logic; // @[Conditional.scala 38:67:@73.18]
  assign _GEN_12 = _T_48 ? _GEN_8 : ack_cpus_ok; // @[Conditional.scala 38:67:@73.18]
  assign _GEN_13 = _T_48 ? _GEN_9 : state; // @[Conditional.scala 38:67:@73.18]
  assign _GEN_14 = _T_43 ? _GEN_4 : _GEN_13; // @[Conditional.scala 38:67:@63.16]
  assign _GEN_15 = _T_43 ? _GEN_5 : _GEN_11; // @[Conditional.scala 38:67:@63.16]
  assign _GEN_16 = _T_43 ? _GEN_6 : _GEN_10; // @[Conditional.scala 38:67:@63.16]
  assign _GEN_17 = _T_43 ? ack_cpus_ok : _GEN_12; // @[Conditional.scala 38:67:@63.16]
  assign _GEN_18 = _T_42 ? _GEN_3 : _GEN_14; // @[Conditional.scala 38:67:@56.14]
  assign _GEN_19 = _T_42 ? reset_routing_logic : _GEN_15; // @[Conditional.scala 38:67:@56.14]
  assign _GEN_20 = _T_42 ? reset_cpus : _GEN_16; // @[Conditional.scala 38:67:@56.14]
  assign _GEN_21 = _T_42 ? ack_cpus_ok : _GEN_17; // @[Conditional.scala 38:67:@56.14]
  assign _GEN_22 = _T_39 ? 3'h5 : _GEN_18; // @[Conditional.scala 38:67:@49.12]
  assign _GEN_23 = _T_39 ? 1'h1 : _GEN_20; // @[Conditional.scala 38:67:@49.12]
  assign _GEN_24 = _T_39 ? 1'h0 : stop_cpus; // @[Conditional.scala 38:67:@49.12]
  assign _GEN_25 = _T_39 ? reset_routing_logic : _GEN_19; // @[Conditional.scala 38:67:@49.12]
  assign _GEN_26 = _T_39 ? ack_cpus_ok : _GEN_21; // @[Conditional.scala 38:67:@49.12]
  assign _GEN_27 = _T_37 ? 3'h4 : _GEN_22; // @[Conditional.scala 38:67:@43.10]
  assign _GEN_28 = _T_37 ? 1'h0 : latch_regs; // @[Conditional.scala 38:67:@43.10]
  assign _GEN_29 = _T_37 ? reset_cpus : _GEN_23; // @[Conditional.scala 38:67:@43.10]
  assign _GEN_30 = _T_37 ? stop_cpus : _GEN_24; // @[Conditional.scala 38:67:@43.10]
  assign _GEN_31 = _T_37 ? reset_routing_logic : _GEN_25; // @[Conditional.scala 38:67:@43.10]
  assign _GEN_32 = _T_37 ? ack_cpus_ok : _GEN_26; // @[Conditional.scala 38:67:@43.10]
  assign _GEN_33 = _T_33 ? _GEN_1 : _GEN_27; // @[Conditional.scala 38:67:@34.8]
  assign _GEN_34 = _T_33 ? _GEN_2 : _GEN_28; // @[Conditional.scala 38:67:@34.8]
  assign _GEN_35 = _T_33 ? reset_cpus : _GEN_29; // @[Conditional.scala 38:67:@34.8]
  assign _GEN_36 = _T_33 ? stop_cpus : _GEN_30; // @[Conditional.scala 38:67:@34.8]
  assign _GEN_37 = _T_33 ? reset_routing_logic : _GEN_31; // @[Conditional.scala 38:67:@34.8]
  assign _GEN_38 = _T_33 ? ack_cpus_ok : _GEN_32; // @[Conditional.scala 38:67:@34.8]
  assign _GEN_39 = _T_30 ? 1'h1 : _GEN_36; // @[Conditional.scala 38:67:@27.6]
  assign _GEN_40 = _T_30 ? 3'h2 : _GEN_33; // @[Conditional.scala 38:67:@27.6]
  assign _GEN_41 = _T_30 ? 1'h1 : reset_to_recovery; // @[Conditional.scala 38:67:@27.6]
  assign _GEN_42 = _T_30 ? latch_regs : _GEN_34; // @[Conditional.scala 38:67:@27.6]
  assign _GEN_43 = _T_30 ? reset_cpus : _GEN_35; // @[Conditional.scala 38:67:@27.6]
  assign _GEN_44 = _T_30 ? reset_routing_logic : _GEN_37; // @[Conditional.scala 38:67:@27.6]
  assign _GEN_45 = _T_30 ? ack_cpus_ok : _GEN_38; // @[Conditional.scala 38:67:@27.6]
  assign _GEN_46 = _T_25 ? 1'h0 : _GEN_39; // @[Conditional.scala 39:58:@16.4]
  assign _GEN_47 = _T_25 ? 1'h0 : _GEN_45; // @[Conditional.scala 39:58:@16.4]
  assign _GEN_48 = _T_25 ? 1'h0 : _GEN_41; // @[Conditional.scala 39:58:@16.4]
  assign _GEN_49 = _T_25 ? 1'h0 : _GEN_44; // @[Conditional.scala 39:58:@16.4]
  assign _GEN_50 = _T_25 ? _GEN_0 : _GEN_40; // @[Conditional.scala 39:58:@16.4]
  assign _GEN_51 = _T_25 ? latch_regs : _GEN_42; // @[Conditional.scala 39:58:@16.4]
  assign _GEN_52 = _T_25 ? reset_cpus : _GEN_43; // @[Conditional.scala 39:58:@16.4]
  assign io_ack_cpus_ok = ack_cpus_ok;
  assign io_stop_cpus = stop_cpus;
  assign io_latch_regs = latch_regs;
  assign io_reset_to_recovery = reset_to_recovery;
  assign io_reset_cpus = reset_cpus;
  assign io_reset_routing_logic = reset_routing_logic;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  state = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  ack_cpus_ok = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  stop_cpus = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  latch_regs = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  reset_to_recovery = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  reset_cpus = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  reset_routing_logic = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 3'h0;
    end else begin
      if (_T_25) begin
        if (io_fault) begin
          state <= 3'h1;
        end
      end else begin
        if (_T_30) begin
          state <= 3'h2;
        end else begin
          if (_T_33) begin
            if (_T_35) begin
              state <= 3'h3;
            end
          end else begin
            if (_T_37) begin
              state <= 3'h4;
            end else begin
              if (_T_39) begin
                state <= 3'h5;
              end else begin
                if (_T_42) begin
                  if (io_reset_pending) begin
                    state <= 3'h6;
                  end
                end else begin
                  if (_T_43) begin
                    if (_T_45) begin
                      state <= 3'h7;
                    end
                  end else begin
                    if (_T_48) begin
                      if (io_cpus_ok) begin
                        state <= 3'h0;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      ack_cpus_ok <= 1'h0;
    end else begin
      if (_T_25) begin
        ack_cpus_ok <= 1'h0;
      end else begin
        if (!(_T_30)) begin
          if (!(_T_33)) begin
            if (!(_T_37)) begin
              if (!(_T_39)) begin
                if (!(_T_42)) begin
                  if (!(_T_43)) begin
                    if (_T_48) begin
                      if (io_cpus_ok) begin
                        ack_cpus_ok <= 1'h1;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      stop_cpus <= 1'h0;
    end else begin
      if (_T_25) begin
        stop_cpus <= 1'h0;
      end else begin
        if (_T_30) begin
          stop_cpus <= 1'h1;
        end else begin
          if (!(_T_33)) begin
            if (!(_T_37)) begin
              if (_T_39) begin
                stop_cpus <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      latch_regs <= 1'h0;
    end else begin
      if (!(_T_25)) begin
        if (!(_T_30)) begin
          if (_T_33) begin
            if (_T_35) begin
              latch_regs <= 1'h1;
            end
          end else begin
            if (_T_37) begin
              latch_regs <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      reset_to_recovery <= 1'h0;
    end else begin
      if (_T_25) begin
        reset_to_recovery <= 1'h0;
      end else begin
        if (_T_30) begin
          reset_to_recovery <= 1'h1;
        end
      end
    end
    if (reset) begin
      reset_cpus <= 1'h0;
    end else begin
      if (!(_T_25)) begin
        if (!(_T_30)) begin
          if (!(_T_33)) begin
            if (!(_T_37)) begin
              if (_T_39) begin
                reset_cpus <= 1'h1;
              end else begin
                if (!(_T_42)) begin
                  if (_T_43) begin
                    if (_T_45) begin
                      reset_cpus <= 1'h0;
                    end
                  end else begin
                    if (_T_48) begin
                      reset_cpus <= 1'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      reset_routing_logic <= 1'h0;
    end else begin
      if (_T_25) begin
        reset_routing_logic <= 1'h0;
      end else begin
        if (!(_T_30)) begin
          if (!(_T_33)) begin
            if (!(_T_37)) begin
              if (!(_T_39)) begin
                if (!(_T_42)) begin
                  if (_T_43) begin
                    if (_T_45) begin
                      reset_routing_logic <= 1'h1;
                    end
                  end else begin
                    if (_T_48) begin
                      if (io_cpus_ok) begin
                        reset_routing_logic <= 1'h0;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module signalHolder( // @[:@88.2]
  input   clock, // @[:@89.4]
  input   io_rst, // @[:@91.4]
  output  io_o, // @[:@91.4]
  input   io_i // @[:@91.4]
);
  reg [6:0] value; // @[Counter.scala 17:33:@93.4]
  reg [31:0] _RAND_0;
  reg  _T_9; // @[FaultDetector.scala 104:23:@94.4]
  reg [31:0] _RAND_1;
  wire  _T_12; // @[Counter.scala 25:24:@97.6]
  wire [7:0] _T_14; // @[Counter.scala 26:22:@98.6]
  wire [6:0] _T_15; // @[Counter.scala 26:22:@99.6]
  wire [6:0] _GEN_0; // @[Counter.scala 28:21:@101.6]
  wire  _GEN_1; // @[FaultDetector.scala 107:25:@104.6]
  wire [6:0] _GEN_2; // @[FaultDetector.scala 106:23:@96.4]
  wire  _GEN_3; // @[FaultDetector.scala 106:23:@96.4]
  wire  _T_18; // @[FaultDetector.scala 111:20:@108.4]
  wire  _T_19; // @[FaultDetector.scala 111:18:@109.4]
  assign _T_12 = value == 7'h63; // @[Counter.scala 25:24:@97.6]
  assign _T_14 = value + 7'h1; // @[Counter.scala 26:22:@98.6]
  assign _T_15 = _T_14[6:0]; // @[Counter.scala 26:22:@99.6]
  assign _GEN_0 = _T_12 ? 7'h0 : _T_15; // @[Counter.scala 28:21:@101.6]
  assign _GEN_1 = _T_12 ? 1'h1 : _T_9; // @[FaultDetector.scala 107:25:@104.6]
  assign _GEN_2 = io_i ? _GEN_0 : value; // @[FaultDetector.scala 106:23:@96.4]
  assign _GEN_3 = io_i ? _GEN_1 : _T_9; // @[FaultDetector.scala 106:23:@96.4]
  assign _T_18 = ~ _T_9; // @[FaultDetector.scala 111:20:@108.4]
  assign _T_19 = io_i & _T_18; // @[FaultDetector.scala 111:18:@109.4]
  assign io_o = _T_19;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  value = _RAND_0[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_9 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (io_rst) begin
      value <= 7'h0;
    end else begin
      if (io_i) begin
        if (_T_12) begin
          value <= 7'h0;
        end else begin
          value <= _T_15;
        end
      end
    end
    if (io_rst) begin
      _T_9 <= 1'h0;
    end else begin
      if (io_i) begin
        if (_T_12) begin
          _T_9 <= 1'h1;
        end
      end
    end
  end
endmodule
module FaultDetector( // @[:@256.2]
  input         clock, // @[:@257.4]
  input         reset, // @[:@258.4]
  output [2:0]  io_invalid, // @[:@259.4]
  output        io_cpu0_axi4_aw_ready, // @[:@259.4]
  input         io_cpu0_axi4_aw_valid, // @[:@259.4]
  input  [3:0]  io_cpu0_axi4_aw_bits_id, // @[:@259.4]
  input  [31:0] io_cpu0_axi4_aw_bits_addr, // @[:@259.4]
  input  [7:0]  io_cpu0_axi4_aw_bits_len, // @[:@259.4]
  input  [2:0]  io_cpu0_axi4_aw_bits_size, // @[:@259.4]
  input  [1:0]  io_cpu0_axi4_aw_bits_burst, // @[:@259.4]
  input         io_cpu0_axi4_aw_bits_lock, // @[:@259.4]
  input  [3:0]  io_cpu0_axi4_aw_bits_cache, // @[:@259.4]
  input  [2:0]  io_cpu0_axi4_aw_bits_prot, // @[:@259.4]
  input  [3:0]  io_cpu0_axi4_aw_bits_qos, // @[:@259.4]
  output        io_cpu0_axi4_w_ready, // @[:@259.4]
  input         io_cpu0_axi4_w_valid, // @[:@259.4]
  input  [31:0] io_cpu0_axi4_w_bits_data, // @[:@259.4]
  input  [3:0]  io_cpu0_axi4_w_bits_strb, // @[:@259.4]
  input         io_cpu0_axi4_w_bits_last, // @[:@259.4]
  input         io_cpu0_axi4_b_ready, // @[:@259.4]
  output        io_cpu0_axi4_b_valid, // @[:@259.4]
  output [3:0]  io_cpu0_axi4_b_bits_id, // @[:@259.4]
  output [1:0]  io_cpu0_axi4_b_bits_resp, // @[:@259.4]
  output        io_cpu0_axi4_ar_ready, // @[:@259.4]
  input         io_cpu0_axi4_ar_valid, // @[:@259.4]
  input  [3:0]  io_cpu0_axi4_ar_bits_id, // @[:@259.4]
  input  [31:0] io_cpu0_axi4_ar_bits_addr, // @[:@259.4]
  input  [7:0]  io_cpu0_axi4_ar_bits_len, // @[:@259.4]
  input  [2:0]  io_cpu0_axi4_ar_bits_size, // @[:@259.4]
  input  [1:0]  io_cpu0_axi4_ar_bits_burst, // @[:@259.4]
  input         io_cpu0_axi4_ar_bits_lock, // @[:@259.4]
  input  [3:0]  io_cpu0_axi4_ar_bits_cache, // @[:@259.4]
  input  [2:0]  io_cpu0_axi4_ar_bits_prot, // @[:@259.4]
  input  [3:0]  io_cpu0_axi4_ar_bits_qos, // @[:@259.4]
  input         io_cpu0_axi4_r_ready, // @[:@259.4]
  output        io_cpu0_axi4_r_valid, // @[:@259.4]
  output [3:0]  io_cpu0_axi4_r_bits_id, // @[:@259.4]
  output [31:0] io_cpu0_axi4_r_bits_data, // @[:@259.4]
  output [1:0]  io_cpu0_axi4_r_bits_resp, // @[:@259.4]
  output        io_cpu0_axi4_r_bits_last, // @[:@259.4]
  output        io_cpu1_axi4_aw_ready, // @[:@259.4]
  input         io_cpu1_axi4_aw_valid, // @[:@259.4]
  input  [3:0]  io_cpu1_axi4_aw_bits_id, // @[:@259.4]
  input  [31:0] io_cpu1_axi4_aw_bits_addr, // @[:@259.4]
  input  [7:0]  io_cpu1_axi4_aw_bits_len, // @[:@259.4]
  input  [2:0]  io_cpu1_axi4_aw_bits_size, // @[:@259.4]
  input  [1:0]  io_cpu1_axi4_aw_bits_burst, // @[:@259.4]
  input         io_cpu1_axi4_aw_bits_lock, // @[:@259.4]
  input  [3:0]  io_cpu1_axi4_aw_bits_cache, // @[:@259.4]
  input  [2:0]  io_cpu1_axi4_aw_bits_prot, // @[:@259.4]
  input  [3:0]  io_cpu1_axi4_aw_bits_qos, // @[:@259.4]
  output        io_cpu1_axi4_w_ready, // @[:@259.4]
  input         io_cpu1_axi4_w_valid, // @[:@259.4]
  input  [31:0] io_cpu1_axi4_w_bits_data, // @[:@259.4]
  input  [3:0]  io_cpu1_axi4_w_bits_strb, // @[:@259.4]
  input         io_cpu1_axi4_w_bits_last, // @[:@259.4]
  input         io_cpu1_axi4_b_ready, // @[:@259.4]
  output        io_cpu1_axi4_b_valid, // @[:@259.4]
  output [3:0]  io_cpu1_axi4_b_bits_id, // @[:@259.4]
  output [1:0]  io_cpu1_axi4_b_bits_resp, // @[:@259.4]
  output        io_cpu1_axi4_ar_ready, // @[:@259.4]
  input         io_cpu1_axi4_ar_valid, // @[:@259.4]
  input  [3:0]  io_cpu1_axi4_ar_bits_id, // @[:@259.4]
  input  [31:0] io_cpu1_axi4_ar_bits_addr, // @[:@259.4]
  input  [7:0]  io_cpu1_axi4_ar_bits_len, // @[:@259.4]
  input  [2:0]  io_cpu1_axi4_ar_bits_size, // @[:@259.4]
  input  [1:0]  io_cpu1_axi4_ar_bits_burst, // @[:@259.4]
  input         io_cpu1_axi4_ar_bits_lock, // @[:@259.4]
  input  [3:0]  io_cpu1_axi4_ar_bits_cache, // @[:@259.4]
  input  [2:0]  io_cpu1_axi4_ar_bits_prot, // @[:@259.4]
  input  [3:0]  io_cpu1_axi4_ar_bits_qos, // @[:@259.4]
  input         io_cpu1_axi4_r_ready, // @[:@259.4]
  output        io_cpu1_axi4_r_valid, // @[:@259.4]
  output [3:0]  io_cpu1_axi4_r_bits_id, // @[:@259.4]
  output [31:0] io_cpu1_axi4_r_bits_data, // @[:@259.4]
  output [1:0]  io_cpu1_axi4_r_bits_resp, // @[:@259.4]
  output        io_cpu1_axi4_r_bits_last, // @[:@259.4]
  output        io_cpu2_axi4_aw_ready, // @[:@259.4]
  input         io_cpu2_axi4_aw_valid, // @[:@259.4]
  input  [3:0]  io_cpu2_axi4_aw_bits_id, // @[:@259.4]
  input  [31:0] io_cpu2_axi4_aw_bits_addr, // @[:@259.4]
  input  [7:0]  io_cpu2_axi4_aw_bits_len, // @[:@259.4]
  input  [2:0]  io_cpu2_axi4_aw_bits_size, // @[:@259.4]
  input  [1:0]  io_cpu2_axi4_aw_bits_burst, // @[:@259.4]
  input         io_cpu2_axi4_aw_bits_lock, // @[:@259.4]
  input  [3:0]  io_cpu2_axi4_aw_bits_cache, // @[:@259.4]
  input  [2:0]  io_cpu2_axi4_aw_bits_prot, // @[:@259.4]
  input  [3:0]  io_cpu2_axi4_aw_bits_qos, // @[:@259.4]
  output        io_cpu2_axi4_w_ready, // @[:@259.4]
  input         io_cpu2_axi4_w_valid, // @[:@259.4]
  input  [31:0] io_cpu2_axi4_w_bits_data, // @[:@259.4]
  input  [3:0]  io_cpu2_axi4_w_bits_strb, // @[:@259.4]
  input         io_cpu2_axi4_w_bits_last, // @[:@259.4]
  input         io_cpu2_axi4_b_ready, // @[:@259.4]
  output        io_cpu2_axi4_b_valid, // @[:@259.4]
  output [3:0]  io_cpu2_axi4_b_bits_id, // @[:@259.4]
  output [1:0]  io_cpu2_axi4_b_bits_resp, // @[:@259.4]
  output        io_cpu2_axi4_ar_ready, // @[:@259.4]
  input         io_cpu2_axi4_ar_valid, // @[:@259.4]
  input  [3:0]  io_cpu2_axi4_ar_bits_id, // @[:@259.4]
  input  [31:0] io_cpu2_axi4_ar_bits_addr, // @[:@259.4]
  input  [7:0]  io_cpu2_axi4_ar_bits_len, // @[:@259.4]
  input  [2:0]  io_cpu2_axi4_ar_bits_size, // @[:@259.4]
  input  [1:0]  io_cpu2_axi4_ar_bits_burst, // @[:@259.4]
  input         io_cpu2_axi4_ar_bits_lock, // @[:@259.4]
  input  [3:0]  io_cpu2_axi4_ar_bits_cache, // @[:@259.4]
  input  [2:0]  io_cpu2_axi4_ar_bits_prot, // @[:@259.4]
  input  [3:0]  io_cpu2_axi4_ar_bits_qos, // @[:@259.4]
  input         io_cpu2_axi4_r_ready, // @[:@259.4]
  output        io_cpu2_axi4_r_valid, // @[:@259.4]
  output [3:0]  io_cpu2_axi4_r_bits_id, // @[:@259.4]
  output [31:0] io_cpu2_axi4_r_bits_data, // @[:@259.4]
  output [1:0]  io_cpu2_axi4_r_bits_resp, // @[:@259.4]
  output        io_cpu2_axi4_r_bits_last, // @[:@259.4]
  input         io_out_axi4_aw_ready, // @[:@259.4]
  output        io_out_axi4_aw_valid, // @[:@259.4]
  output [3:0]  io_out_axi4_aw_bits_id, // @[:@259.4]
  output [31:0] io_out_axi4_aw_bits_addr, // @[:@259.4]
  output [7:0]  io_out_axi4_aw_bits_len, // @[:@259.4]
  output [2:0]  io_out_axi4_aw_bits_size, // @[:@259.4]
  output [1:0]  io_out_axi4_aw_bits_burst, // @[:@259.4]
  output        io_out_axi4_aw_bits_lock, // @[:@259.4]
  output [3:0]  io_out_axi4_aw_bits_cache, // @[:@259.4]
  output [2:0]  io_out_axi4_aw_bits_prot, // @[:@259.4]
  output [3:0]  io_out_axi4_aw_bits_qos, // @[:@259.4]
  input         io_out_axi4_w_ready, // @[:@259.4]
  output        io_out_axi4_w_valid, // @[:@259.4]
  output [31:0] io_out_axi4_w_bits_data, // @[:@259.4]
  output [3:0]  io_out_axi4_w_bits_strb, // @[:@259.4]
  output        io_out_axi4_w_bits_last, // @[:@259.4]
  output        io_out_axi4_b_ready, // @[:@259.4]
  input         io_out_axi4_b_valid, // @[:@259.4]
  input  [3:0]  io_out_axi4_b_bits_id, // @[:@259.4]
  input  [1:0]  io_out_axi4_b_bits_resp, // @[:@259.4]
  input         io_out_axi4_ar_ready, // @[:@259.4]
  output        io_out_axi4_ar_valid, // @[:@259.4]
  output [3:0]  io_out_axi4_ar_bits_id, // @[:@259.4]
  output [31:0] io_out_axi4_ar_bits_addr, // @[:@259.4]
  output [7:0]  io_out_axi4_ar_bits_len, // @[:@259.4]
  output [2:0]  io_out_axi4_ar_bits_size, // @[:@259.4]
  output [1:0]  io_out_axi4_ar_bits_burst, // @[:@259.4]
  output        io_out_axi4_ar_bits_lock, // @[:@259.4]
  output [3:0]  io_out_axi4_ar_bits_cache, // @[:@259.4]
  output [2:0]  io_out_axi4_ar_bits_prot, // @[:@259.4]
  output [3:0]  io_out_axi4_ar_bits_qos, // @[:@259.4]
  output        io_out_axi4_r_ready, // @[:@259.4]
  input         io_out_axi4_r_valid, // @[:@259.4]
  input  [3:0]  io_out_axi4_r_bits_id, // @[:@259.4]
  input  [31:0] io_out_axi4_r_bits_data, // @[:@259.4]
  input  [1:0]  io_out_axi4_r_bits_resp, // @[:@259.4]
  input         io_out_axi4_r_bits_last, // @[:@259.4]
  output [2:0]  io_fault_reset_vector, // @[:@259.4]
  output [2:0]  io_reset_cpu, // @[:@259.4]
  output        io_stop_all_cpus, // @[:@259.4]
  output        io_latch_registers, // @[:@259.4]
  output        io_reset_to_recovery, // @[:@259.4]
  input         io_cpu_reset_feedback, // @[:@259.4]
  input         io_disable_reset, // @[:@259.4]
  input  [2:0]  io_reset_routing_logic, // @[:@259.4]
  output        io_cpu_back_online, // @[:@259.4]
  input         io_ack_back_online, // @[:@259.4]
  input         io_cpu_in_interrupt // @[:@259.4]
);
  wire  cpu_repair_clock; // @[FaultDetector.scala 394:26:@261.4]
  wire  cpu_repair_reset; // @[FaultDetector.scala 394:26:@261.4]
  wire  cpu_repair_io_fault; // @[FaultDetector.scala 394:26:@261.4]
  wire  cpu_repair_io_cpus_ok; // @[FaultDetector.scala 394:26:@261.4]
  wire  cpu_repair_io_reset_pending; // @[FaultDetector.scala 394:26:@261.4]
  wire  cpu_repair_io_ack_cpus_ok; // @[FaultDetector.scala 394:26:@261.4]
  wire  cpu_repair_io_stop_cpus; // @[FaultDetector.scala 394:26:@261.4]
  wire  cpu_repair_io_latch_regs; // @[FaultDetector.scala 394:26:@261.4]
  wire  cpu_repair_io_reset_to_recovery; // @[FaultDetector.scala 394:26:@261.4]
  wire  cpu_repair_io_reset_cpus; // @[FaultDetector.scala 394:26:@261.4]
  wire  cpu_repair_io_reset_routing_logic; // @[FaultDetector.scala 394:26:@261.4]
  wire  cpu_repair_io_cpu_in_interrupt; // @[FaultDetector.scala 394:26:@261.4]
  wire  axiBusInternal0_aw_ready; // @[FaultDetector.scala 396:29:@264.4]
  wire  axiBusInternal0_aw_valid; // @[FaultDetector.scala 396:29:@264.4]
  wire [3:0] axiBusInternal0_aw_bits_id; // @[FaultDetector.scala 396:29:@264.4]
  wire [31:0] axiBusInternal0_aw_bits_addr; // @[FaultDetector.scala 396:29:@264.4]
  wire [7:0] axiBusInternal0_aw_bits_len; // @[FaultDetector.scala 396:29:@264.4]
  wire [2:0] axiBusInternal0_aw_bits_size; // @[FaultDetector.scala 396:29:@264.4]
  wire [1:0] axiBusInternal0_aw_bits_burst; // @[FaultDetector.scala 396:29:@264.4]
  wire  axiBusInternal0_aw_bits_lock; // @[FaultDetector.scala 396:29:@264.4]
  wire [3:0] axiBusInternal0_aw_bits_cache; // @[FaultDetector.scala 396:29:@264.4]
  wire [2:0] axiBusInternal0_aw_bits_prot; // @[FaultDetector.scala 396:29:@264.4]
  wire [3:0] axiBusInternal0_aw_bits_qos; // @[FaultDetector.scala 396:29:@264.4]
  wire  axiBusInternal0_w_ready; // @[FaultDetector.scala 396:29:@264.4]
  wire  axiBusInternal0_w_valid; // @[FaultDetector.scala 396:29:@264.4]
  wire [31:0] axiBusInternal0_w_bits_data; // @[FaultDetector.scala 396:29:@264.4]
  wire [3:0] axiBusInternal0_w_bits_strb; // @[FaultDetector.scala 396:29:@264.4]
  wire  axiBusInternal0_w_bits_last; // @[FaultDetector.scala 396:29:@264.4]
  wire  axiBusInternal0_b_ready; // @[FaultDetector.scala 396:29:@264.4]
  wire  axiBusInternal0_b_valid; // @[FaultDetector.scala 396:29:@264.4]
  wire [3:0] axiBusInternal0_b_bits_id; // @[FaultDetector.scala 396:29:@264.4]
  wire [1:0] axiBusInternal0_b_bits_resp; // @[FaultDetector.scala 396:29:@264.4]
  wire  axiBusInternal0_ar_ready; // @[FaultDetector.scala 396:29:@264.4]
  wire  axiBusInternal0_ar_valid; // @[FaultDetector.scala 396:29:@264.4]
  wire [3:0] axiBusInternal0_ar_bits_id; // @[FaultDetector.scala 396:29:@264.4]
  wire [31:0] axiBusInternal0_ar_bits_addr; // @[FaultDetector.scala 396:29:@264.4]
  wire [7:0] axiBusInternal0_ar_bits_len; // @[FaultDetector.scala 396:29:@264.4]
  wire [2:0] axiBusInternal0_ar_bits_size; // @[FaultDetector.scala 396:29:@264.4]
  wire [1:0] axiBusInternal0_ar_bits_burst; // @[FaultDetector.scala 396:29:@264.4]
  wire  axiBusInternal0_ar_bits_lock; // @[FaultDetector.scala 396:29:@264.4]
  wire [3:0] axiBusInternal0_ar_bits_cache; // @[FaultDetector.scala 396:29:@264.4]
  wire [2:0] axiBusInternal0_ar_bits_prot; // @[FaultDetector.scala 396:29:@264.4]
  wire [3:0] axiBusInternal0_ar_bits_qos; // @[FaultDetector.scala 396:29:@264.4]
  wire  axiBusInternal0_r_ready; // @[FaultDetector.scala 396:29:@264.4]
  wire  axiBusInternal0_r_valid; // @[FaultDetector.scala 396:29:@264.4]
  wire [3:0] axiBusInternal0_r_bits_id; // @[FaultDetector.scala 396:29:@264.4]
  wire [31:0] axiBusInternal0_r_bits_data; // @[FaultDetector.scala 396:29:@264.4]
  wire [1:0] axiBusInternal0_r_bits_resp; // @[FaultDetector.scala 396:29:@264.4]
  wire  axiBusInternal0_r_bits_last; // @[FaultDetector.scala 396:29:@264.4]
  wire  axiBusInternal1_aw_ready; // @[FaultDetector.scala 397:29:@265.4]
  wire  axiBusInternal1_aw_valid; // @[FaultDetector.scala 397:29:@265.4]
  wire [3:0] axiBusInternal1_aw_bits_id; // @[FaultDetector.scala 397:29:@265.4]
  wire [31:0] axiBusInternal1_aw_bits_addr; // @[FaultDetector.scala 397:29:@265.4]
  wire [7:0] axiBusInternal1_aw_bits_len; // @[FaultDetector.scala 397:29:@265.4]
  wire [2:0] axiBusInternal1_aw_bits_size; // @[FaultDetector.scala 397:29:@265.4]
  wire [1:0] axiBusInternal1_aw_bits_burst; // @[FaultDetector.scala 397:29:@265.4]
  wire  axiBusInternal1_aw_bits_lock; // @[FaultDetector.scala 397:29:@265.4]
  wire [3:0] axiBusInternal1_aw_bits_cache; // @[FaultDetector.scala 397:29:@265.4]
  wire [2:0] axiBusInternal1_aw_bits_prot; // @[FaultDetector.scala 397:29:@265.4]
  wire [3:0] axiBusInternal1_aw_bits_qos; // @[FaultDetector.scala 397:29:@265.4]
  wire  axiBusInternal1_w_ready; // @[FaultDetector.scala 397:29:@265.4]
  wire  axiBusInternal1_w_valid; // @[FaultDetector.scala 397:29:@265.4]
  wire [31:0] axiBusInternal1_w_bits_data; // @[FaultDetector.scala 397:29:@265.4]
  wire [3:0] axiBusInternal1_w_bits_strb; // @[FaultDetector.scala 397:29:@265.4]
  wire  axiBusInternal1_w_bits_last; // @[FaultDetector.scala 397:29:@265.4]
  wire  axiBusInternal1_b_ready; // @[FaultDetector.scala 397:29:@265.4]
  wire  axiBusInternal1_b_valid; // @[FaultDetector.scala 397:29:@265.4]
  wire [3:0] axiBusInternal1_b_bits_id; // @[FaultDetector.scala 397:29:@265.4]
  wire [1:0] axiBusInternal1_b_bits_resp; // @[FaultDetector.scala 397:29:@265.4]
  wire  axiBusInternal1_ar_ready; // @[FaultDetector.scala 397:29:@265.4]
  wire  axiBusInternal1_ar_valid; // @[FaultDetector.scala 397:29:@265.4]
  wire [3:0] axiBusInternal1_ar_bits_id; // @[FaultDetector.scala 397:29:@265.4]
  wire [31:0] axiBusInternal1_ar_bits_addr; // @[FaultDetector.scala 397:29:@265.4]
  wire [7:0] axiBusInternal1_ar_bits_len; // @[FaultDetector.scala 397:29:@265.4]
  wire [2:0] axiBusInternal1_ar_bits_size; // @[FaultDetector.scala 397:29:@265.4]
  wire [1:0] axiBusInternal1_ar_bits_burst; // @[FaultDetector.scala 397:29:@265.4]
  wire  axiBusInternal1_ar_bits_lock; // @[FaultDetector.scala 397:29:@265.4]
  wire [3:0] axiBusInternal1_ar_bits_cache; // @[FaultDetector.scala 397:29:@265.4]
  wire [2:0] axiBusInternal1_ar_bits_prot; // @[FaultDetector.scala 397:29:@265.4]
  wire [3:0] axiBusInternal1_ar_bits_qos; // @[FaultDetector.scala 397:29:@265.4]
  wire  axiBusInternal1_r_ready; // @[FaultDetector.scala 397:29:@265.4]
  wire  axiBusInternal1_r_valid; // @[FaultDetector.scala 397:29:@265.4]
  wire [3:0] axiBusInternal1_r_bits_id; // @[FaultDetector.scala 397:29:@265.4]
  wire [31:0] axiBusInternal1_r_bits_data; // @[FaultDetector.scala 397:29:@265.4]
  wire [1:0] axiBusInternal1_r_bits_resp; // @[FaultDetector.scala 397:29:@265.4]
  wire  axiBusInternal1_r_bits_last; // @[FaultDetector.scala 397:29:@265.4]
  wire  axiBusInternal2_aw_ready; // @[FaultDetector.scala 398:29:@266.4]
  wire  axiBusInternal2_aw_valid; // @[FaultDetector.scala 398:29:@266.4]
  wire [3:0] axiBusInternal2_aw_bits_id; // @[FaultDetector.scala 398:29:@266.4]
  wire [31:0] axiBusInternal2_aw_bits_addr; // @[FaultDetector.scala 398:29:@266.4]
  wire [7:0] axiBusInternal2_aw_bits_len; // @[FaultDetector.scala 398:29:@266.4]
  wire [2:0] axiBusInternal2_aw_bits_size; // @[FaultDetector.scala 398:29:@266.4]
  wire [1:0] axiBusInternal2_aw_bits_burst; // @[FaultDetector.scala 398:29:@266.4]
  wire  axiBusInternal2_aw_bits_lock; // @[FaultDetector.scala 398:29:@266.4]
  wire [3:0] axiBusInternal2_aw_bits_cache; // @[FaultDetector.scala 398:29:@266.4]
  wire [2:0] axiBusInternal2_aw_bits_prot; // @[FaultDetector.scala 398:29:@266.4]
  wire [3:0] axiBusInternal2_aw_bits_qos; // @[FaultDetector.scala 398:29:@266.4]
  wire  axiBusInternal2_w_ready; // @[FaultDetector.scala 398:29:@266.4]
  wire  axiBusInternal2_w_valid; // @[FaultDetector.scala 398:29:@266.4]
  wire [31:0] axiBusInternal2_w_bits_data; // @[FaultDetector.scala 398:29:@266.4]
  wire [3:0] axiBusInternal2_w_bits_strb; // @[FaultDetector.scala 398:29:@266.4]
  wire  axiBusInternal2_w_bits_last; // @[FaultDetector.scala 398:29:@266.4]
  wire  axiBusInternal2_b_ready; // @[FaultDetector.scala 398:29:@266.4]
  wire  axiBusInternal2_b_valid; // @[FaultDetector.scala 398:29:@266.4]
  wire [3:0] axiBusInternal2_b_bits_id; // @[FaultDetector.scala 398:29:@266.4]
  wire [1:0] axiBusInternal2_b_bits_resp; // @[FaultDetector.scala 398:29:@266.4]
  wire  axiBusInternal2_ar_ready; // @[FaultDetector.scala 398:29:@266.4]
  wire  axiBusInternal2_ar_valid; // @[FaultDetector.scala 398:29:@266.4]
  wire [3:0] axiBusInternal2_ar_bits_id; // @[FaultDetector.scala 398:29:@266.4]
  wire [31:0] axiBusInternal2_ar_bits_addr; // @[FaultDetector.scala 398:29:@266.4]
  wire [7:0] axiBusInternal2_ar_bits_len; // @[FaultDetector.scala 398:29:@266.4]
  wire [2:0] axiBusInternal2_ar_bits_size; // @[FaultDetector.scala 398:29:@266.4]
  wire [1:0] axiBusInternal2_ar_bits_burst; // @[FaultDetector.scala 398:29:@266.4]
  wire  axiBusInternal2_ar_bits_lock; // @[FaultDetector.scala 398:29:@266.4]
  wire [3:0] axiBusInternal2_ar_bits_cache; // @[FaultDetector.scala 398:29:@266.4]
  wire [2:0] axiBusInternal2_ar_bits_prot; // @[FaultDetector.scala 398:29:@266.4]
  wire [3:0] axiBusInternal2_ar_bits_qos; // @[FaultDetector.scala 398:29:@266.4]
  wire  axiBusInternal2_r_ready; // @[FaultDetector.scala 398:29:@266.4]
  wire  axiBusInternal2_r_valid; // @[FaultDetector.scala 398:29:@266.4]
  wire [3:0] axiBusInternal2_r_bits_id; // @[FaultDetector.scala 398:29:@266.4]
  wire [31:0] axiBusInternal2_r_bits_data; // @[FaultDetector.scala 398:29:@266.4]
  wire [1:0] axiBusInternal2_r_bits_resp; // @[FaultDetector.scala 398:29:@266.4]
  wire  axiBusInternal2_r_bits_last; // @[FaultDetector.scala 398:29:@266.4]
  wire  reset_logic; // @[FaultDetector.scala 404:25:@267.4]
  wire  reset_routing_0; // @[FaultDetector.scala 405:26:@272.4]
  wire  reset_routing_1; // @[FaultDetector.scala 405:26:@272.4]
  wire  reset_routing_2; // @[FaultDetector.scala 405:26:@272.4]
  wire  logic_reset_hold_0_clock; // @[FaultDetector.scala 406:50:@276.4]
  wire  logic_reset_hold_0_io_rst; // @[FaultDetector.scala 406:50:@276.4]
  wire  logic_reset_hold_0_io_o; // @[FaultDetector.scala 406:50:@276.4]
  wire  logic_reset_hold_0_io_i; // @[FaultDetector.scala 406:50:@276.4]
  wire  logic_reset_hold_1_clock; // @[FaultDetector.scala 406:87:@279.4]
  wire  logic_reset_hold_1_io_rst; // @[FaultDetector.scala 406:87:@279.4]
  wire  logic_reset_hold_1_io_o; // @[FaultDetector.scala 406:87:@279.4]
  wire  logic_reset_hold_1_io_i; // @[FaultDetector.scala 406:87:@279.4]
  wire  logic_reset_hold_2_clock; // @[FaultDetector.scala 406:124:@282.4]
  wire  logic_reset_hold_2_io_rst; // @[FaultDetector.scala 406:124:@282.4]
  wire  logic_reset_hold_2_io_o; // @[FaultDetector.scala 406:124:@282.4]
  wire  logic_reset_hold_2_io_i; // @[FaultDetector.scala 406:124:@282.4]
  wire  _T_397; // @[FaultDetector.scala 410:18:@286.4]
  reg  _T_429_aw_ready; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_0;
  reg  _T_429_aw_valid; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_1;
  reg [3:0] _T_429_aw_bits_id; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_2;
  reg [31:0] _T_429_aw_bits_addr; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_3;
  reg [7:0] _T_429_aw_bits_len; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_4;
  reg [2:0] _T_429_aw_bits_size; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_5;
  reg [1:0] _T_429_aw_bits_burst; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_6;
  reg  _T_429_aw_bits_lock; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_7;
  reg [3:0] _T_429_aw_bits_cache; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_8;
  reg [2:0] _T_429_aw_bits_prot; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_9;
  reg [3:0] _T_429_aw_bits_qos; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_10;
  reg  _T_429_w_ready; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_11;
  reg  _T_429_w_valid; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_12;
  reg [31:0] _T_429_w_bits_data; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_13;
  reg [3:0] _T_429_w_bits_strb; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_14;
  reg  _T_429_w_bits_last; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_15;
  reg  _T_429_b_ready; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_16;
  reg  _T_429_b_valid; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_17;
  reg [3:0] _T_429_b_bits_id; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_18;
  reg [1:0] _T_429_b_bits_resp; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_19;
  reg  _T_429_ar_ready; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_20;
  reg  _T_429_ar_valid; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_21;
  reg [3:0] _T_429_ar_bits_id; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_22;
  reg [31:0] _T_429_ar_bits_addr; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_23;
  reg [7:0] _T_429_ar_bits_len; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_24;
  reg [2:0] _T_429_ar_bits_size; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_25;
  reg [1:0] _T_429_ar_bits_burst; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_26;
  reg  _T_429_ar_bits_lock; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_27;
  reg [3:0] _T_429_ar_bits_cache; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_28;
  reg [2:0] _T_429_ar_bits_prot; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_29;
  reg [3:0] _T_429_ar_bits_qos; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_30;
  reg  _T_429_r_ready; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_31;
  reg  _T_429_r_valid; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_32;
  reg [3:0] _T_429_r_bits_id; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_33;
  reg [31:0] _T_429_r_bits_data; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_34;
  reg [1:0] _T_429_r_bits_resp; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_35;
  reg  _T_429_r_bits_last; // @[FaultDetector.scala 117:19:@297.4]
  reg [31:0] _RAND_36;
  reg  _T_487_aw_ready; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_37;
  reg  _T_487_aw_valid; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_38;
  reg [3:0] _T_487_aw_bits_id; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_39;
  reg [31:0] _T_487_aw_bits_addr; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_40;
  reg [7:0] _T_487_aw_bits_len; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_41;
  reg [2:0] _T_487_aw_bits_size; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_42;
  reg [1:0] _T_487_aw_bits_burst; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_43;
  reg  _T_487_aw_bits_lock; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_44;
  reg [3:0] _T_487_aw_bits_cache; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_45;
  reg [2:0] _T_487_aw_bits_prot; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_46;
  reg [3:0] _T_487_aw_bits_qos; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_47;
  reg  _T_487_w_ready; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_48;
  reg  _T_487_w_valid; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_49;
  reg [31:0] _T_487_w_bits_data; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_50;
  reg [3:0] _T_487_w_bits_strb; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_51;
  reg  _T_487_w_bits_last; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_52;
  reg  _T_487_b_ready; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_53;
  reg  _T_487_b_valid; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_54;
  reg [3:0] _T_487_b_bits_id; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_55;
  reg [1:0] _T_487_b_bits_resp; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_56;
  reg  _T_487_ar_ready; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_57;
  reg  _T_487_ar_valid; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_58;
  reg [3:0] _T_487_ar_bits_id; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_59;
  reg [31:0] _T_487_ar_bits_addr; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_60;
  reg [7:0] _T_487_ar_bits_len; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_61;
  reg [2:0] _T_487_ar_bits_size; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_62;
  reg [1:0] _T_487_ar_bits_burst; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_63;
  reg  _T_487_ar_bits_lock; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_64;
  reg [3:0] _T_487_ar_bits_cache; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_65;
  reg [2:0] _T_487_ar_bits_prot; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_66;
  reg [3:0] _T_487_ar_bits_qos; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_67;
  reg  _T_487_r_ready; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_68;
  reg  _T_487_r_valid; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_69;
  reg [3:0] _T_487_r_bits_id; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_70;
  reg [31:0] _T_487_r_bits_data; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_71;
  reg [1:0] _T_487_r_bits_resp; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_72;
  reg  _T_487_r_bits_last; // @[FaultDetector.scala 118:21:@298.4]
  reg [31:0] _RAND_73;
  reg  _T_545_aw_ready; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_74;
  reg  _T_545_aw_valid; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_75;
  reg [3:0] _T_545_aw_bits_id; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_76;
  reg [31:0] _T_545_aw_bits_addr; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_77;
  reg [7:0] _T_545_aw_bits_len; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_78;
  reg [2:0] _T_545_aw_bits_size; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_79;
  reg [1:0] _T_545_aw_bits_burst; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_80;
  reg  _T_545_aw_bits_lock; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_81;
  reg [3:0] _T_545_aw_bits_cache; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_82;
  reg [2:0] _T_545_aw_bits_prot; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_83;
  reg [3:0] _T_545_aw_bits_qos; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_84;
  reg  _T_545_w_ready; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_85;
  reg  _T_545_w_valid; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_86;
  reg [31:0] _T_545_w_bits_data; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_87;
  reg [3:0] _T_545_w_bits_strb; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_88;
  reg  _T_545_w_bits_last; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_89;
  reg  _T_545_b_ready; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_90;
  reg  _T_545_b_valid; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_91;
  reg [3:0] _T_545_b_bits_id; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_92;
  reg [1:0] _T_545_b_bits_resp; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_93;
  reg  _T_545_ar_ready; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_94;
  reg  _T_545_ar_valid; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_95;
  reg [3:0] _T_545_ar_bits_id; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_96;
  reg [31:0] _T_545_ar_bits_addr; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_97;
  reg [7:0] _T_545_ar_bits_len; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_98;
  reg [2:0] _T_545_ar_bits_size; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_99;
  reg [1:0] _T_545_ar_bits_burst; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_100;
  reg  _T_545_ar_bits_lock; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_101;
  reg [3:0] _T_545_ar_bits_cache; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_102;
  reg [2:0] _T_545_ar_bits_prot; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_103;
  reg [3:0] _T_545_ar_bits_qos; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_104;
  reg  _T_545_r_ready; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_105;
  reg  _T_545_r_valid; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_106;
  reg [3:0] _T_545_r_bits_id; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_107;
  reg [31:0] _T_545_r_bits_data; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_108;
  reg [1:0] _T_545_r_bits_resp; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_109;
  reg  _T_545_r_bits_last; // @[FaultDetector.scala 117:19:@299.4]
  reg [31:0] _RAND_110;
  reg  _T_603_aw_ready; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_111;
  reg  _T_603_aw_valid; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_112;
  reg [3:0] _T_603_aw_bits_id; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_113;
  reg [31:0] _T_603_aw_bits_addr; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_114;
  reg [7:0] _T_603_aw_bits_len; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_115;
  reg [2:0] _T_603_aw_bits_size; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_116;
  reg [1:0] _T_603_aw_bits_burst; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_117;
  reg  _T_603_aw_bits_lock; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_118;
  reg [3:0] _T_603_aw_bits_cache; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_119;
  reg [2:0] _T_603_aw_bits_prot; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_120;
  reg [3:0] _T_603_aw_bits_qos; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_121;
  reg  _T_603_w_ready; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_122;
  reg  _T_603_w_valid; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_123;
  reg [31:0] _T_603_w_bits_data; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_124;
  reg [3:0] _T_603_w_bits_strb; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_125;
  reg  _T_603_w_bits_last; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_126;
  reg  _T_603_b_ready; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_127;
  reg  _T_603_b_valid; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_128;
  reg [3:0] _T_603_b_bits_id; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_129;
  reg [1:0] _T_603_b_bits_resp; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_130;
  reg  _T_603_ar_ready; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_131;
  reg  _T_603_ar_valid; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_132;
  reg [3:0] _T_603_ar_bits_id; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_133;
  reg [31:0] _T_603_ar_bits_addr; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_134;
  reg [7:0] _T_603_ar_bits_len; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_135;
  reg [2:0] _T_603_ar_bits_size; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_136;
  reg [1:0] _T_603_ar_bits_burst; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_137;
  reg  _T_603_ar_bits_lock; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_138;
  reg [3:0] _T_603_ar_bits_cache; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_139;
  reg [2:0] _T_603_ar_bits_prot; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_140;
  reg [3:0] _T_603_ar_bits_qos; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_141;
  reg  _T_603_r_ready; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_142;
  reg  _T_603_r_valid; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_143;
  reg [3:0] _T_603_r_bits_id; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_144;
  reg [31:0] _T_603_r_bits_data; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_145;
  reg [1:0] _T_603_r_bits_resp; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_146;
  reg  _T_603_r_bits_last; // @[FaultDetector.scala 118:21:@300.4]
  reg [31:0] _RAND_147;
  reg  _T_661_aw_ready; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_148;
  reg  _T_661_aw_valid; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_149;
  reg [3:0] _T_661_aw_bits_id; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_150;
  reg [31:0] _T_661_aw_bits_addr; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_151;
  reg [7:0] _T_661_aw_bits_len; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_152;
  reg [2:0] _T_661_aw_bits_size; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_153;
  reg [1:0] _T_661_aw_bits_burst; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_154;
  reg  _T_661_aw_bits_lock; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_155;
  reg [3:0] _T_661_aw_bits_cache; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_156;
  reg [2:0] _T_661_aw_bits_prot; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_157;
  reg [3:0] _T_661_aw_bits_qos; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_158;
  reg  _T_661_w_ready; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_159;
  reg  _T_661_w_valid; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_160;
  reg [31:0] _T_661_w_bits_data; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_161;
  reg [3:0] _T_661_w_bits_strb; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_162;
  reg  _T_661_w_bits_last; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_163;
  reg  _T_661_b_ready; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_164;
  reg  _T_661_b_valid; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_165;
  reg [3:0] _T_661_b_bits_id; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_166;
  reg [1:0] _T_661_b_bits_resp; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_167;
  reg  _T_661_ar_ready; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_168;
  reg  _T_661_ar_valid; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_169;
  reg [3:0] _T_661_ar_bits_id; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_170;
  reg [31:0] _T_661_ar_bits_addr; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_171;
  reg [7:0] _T_661_ar_bits_len; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_172;
  reg [2:0] _T_661_ar_bits_size; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_173;
  reg [1:0] _T_661_ar_bits_burst; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_174;
  reg  _T_661_ar_bits_lock; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_175;
  reg [3:0] _T_661_ar_bits_cache; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_176;
  reg [2:0] _T_661_ar_bits_prot; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_177;
  reg [3:0] _T_661_ar_bits_qos; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_178;
  reg  _T_661_r_ready; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_179;
  reg  _T_661_r_valid; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_180;
  reg [3:0] _T_661_r_bits_id; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_181;
  reg [31:0] _T_661_r_bits_data; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_182;
  reg [1:0] _T_661_r_bits_resp; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_183;
  reg  _T_661_r_bits_last; // @[FaultDetector.scala 117:19:@301.4]
  reg [31:0] _RAND_184;
  reg  _T_719_aw_ready; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_185;
  reg  _T_719_aw_valid; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_186;
  reg [3:0] _T_719_aw_bits_id; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_187;
  reg [31:0] _T_719_aw_bits_addr; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_188;
  reg [7:0] _T_719_aw_bits_len; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_189;
  reg [2:0] _T_719_aw_bits_size; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_190;
  reg [1:0] _T_719_aw_bits_burst; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_191;
  reg  _T_719_aw_bits_lock; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_192;
  reg [3:0] _T_719_aw_bits_cache; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_193;
  reg [2:0] _T_719_aw_bits_prot; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_194;
  reg [3:0] _T_719_aw_bits_qos; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_195;
  reg  _T_719_w_ready; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_196;
  reg  _T_719_w_valid; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_197;
  reg [31:0] _T_719_w_bits_data; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_198;
  reg [3:0] _T_719_w_bits_strb; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_199;
  reg  _T_719_w_bits_last; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_200;
  reg  _T_719_b_ready; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_201;
  reg  _T_719_b_valid; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_202;
  reg [3:0] _T_719_b_bits_id; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_203;
  reg [1:0] _T_719_b_bits_resp; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_204;
  reg  _T_719_ar_ready; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_205;
  reg  _T_719_ar_valid; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_206;
  reg [3:0] _T_719_ar_bits_id; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_207;
  reg [31:0] _T_719_ar_bits_addr; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_208;
  reg [7:0] _T_719_ar_bits_len; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_209;
  reg [2:0] _T_719_ar_bits_size; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_210;
  reg [1:0] _T_719_ar_bits_burst; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_211;
  reg  _T_719_ar_bits_lock; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_212;
  reg [3:0] _T_719_ar_bits_cache; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_213;
  reg [2:0] _T_719_ar_bits_prot; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_214;
  reg [3:0] _T_719_ar_bits_qos; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_215;
  reg  _T_719_r_ready; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_216;
  reg  _T_719_r_valid; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_217;
  reg [3:0] _T_719_r_bits_id; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_218;
  reg [31:0] _T_719_r_bits_data; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_219;
  reg [1:0] _T_719_r_bits_resp; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_220;
  reg  _T_719_r_bits_last; // @[FaultDetector.scala 118:21:@302.4]
  reg [31:0] _RAND_221;
  wire  cpu_reset_hold_0_clock; // @[FaultDetector.scala 420:48:@303.4]
  wire  cpu_reset_hold_0_io_rst; // @[FaultDetector.scala 420:48:@303.4]
  wire  cpu_reset_hold_0_io_o; // @[FaultDetector.scala 420:48:@303.4]
  wire  cpu_reset_hold_0_io_i; // @[FaultDetector.scala 420:48:@303.4]
  wire  cpu_reset_hold_1_clock; // @[FaultDetector.scala 420:85:@306.4]
  wire  cpu_reset_hold_1_io_rst; // @[FaultDetector.scala 420:85:@306.4]
  wire  cpu_reset_hold_1_io_o; // @[FaultDetector.scala 420:85:@306.4]
  wire  cpu_reset_hold_1_io_i; // @[FaultDetector.scala 420:85:@306.4]
  wire  cpu_reset_hold_2_clock; // @[FaultDetector.scala 420:122:@309.4]
  wire  cpu_reset_hold_2_io_rst; // @[FaultDetector.scala 420:122:@309.4]
  wire  cpu_reset_hold_2_io_o; // @[FaultDetector.scala 420:122:@309.4]
  wire  cpu_reset_hold_2_io_i; // @[FaultDetector.scala 420:122:@309.4]
  reg [2:0] cpu_reset_im; // @[FaultDetector.scala 421:25:@312.4]
  reg [31:0] _RAND_222;
  wire  cpu_reset_out_0; // @[FaultDetector.scala 423:26:@317.4]
  wire  cpu_reset_out_1; // @[FaultDetector.scala 423:26:@317.4]
  wire  cpu_reset_out_2; // @[FaultDetector.scala 423:26:@317.4]
  wire [1:0] _T_761; // @[FaultDetector.scala 425:52:@321.4]
  wire [2:0] _T_762; // @[FaultDetector.scala 425:52:@322.4]
  wire  _T_764; // @[FaultDetector.scala 425:59:@323.4]
  wire  _T_768_0; // @[FaultDetector.scala 316:25:@324.4]
  wire  _T_768_1; // @[FaultDetector.scala 316:25:@324.4]
  wire  _T_768_2; // @[FaultDetector.scala 316:25:@324.4]
  wire  _T_891_0_0; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_1; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_2; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_3; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_4; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_5; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_6; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_7; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_8; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_9; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_10; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_11; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_12; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_13; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_14; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_15; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_16; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_17; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_18; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_19; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_20; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_21; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_22; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_23; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_24; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_0_25; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_0; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_1; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_2; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_3; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_4; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_5; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_6; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_7; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_8; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_9; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_10; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_11; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_12; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_13; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_14; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_15; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_16; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_17; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_18; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_19; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_20; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_21; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_22; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_23; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_24; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_1_25; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_0; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_1; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_2; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_3; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_4; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_5; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_6; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_7; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_8; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_9; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_10; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_11; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_12; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_13; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_14; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_15; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_16; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_17; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_18; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_19; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_20; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_21; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_22; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_23; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_24; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_891_2_25; // @[FaultDetector.scala 318:29:@325.4]
  wire  _T_1229; // @[FaultDetector.scala 323:43:@326.4]
  wire  _T_1230; // @[FaultDetector.scala 324:42:@328.4]
  wire  _T_1231; // @[FaultDetector.scala 325:43:@330.4]
  wire  _T_1232; // @[FaultDetector.scala 327:42:@332.4]
  wire  _T_1233; // @[FaultDetector.scala 328:42:@334.4]
  wire [3:0] _T_1234; // @[FaultDetector.scala 330:46:@336.4]
  wire  _T_1236; // @[FaultDetector.scala 330:67:@337.4]
  wire [31:0] _T_1237; // @[FaultDetector.scala 331:48:@339.4]
  wire  _T_1239; // @[FaultDetector.scala 331:71:@340.4]
  wire [7:0] _T_1240; // @[FaultDetector.scala 332:47:@342.4]
  wire  _T_1242; // @[FaultDetector.scala 332:69:@343.4]
  wire [2:0] _T_1243; // @[FaultDetector.scala 333:48:@345.4]
  wire  _T_1245; // @[FaultDetector.scala 333:71:@346.4]
  wire [1:0] _T_1246; // @[FaultDetector.scala 334:49:@348.4]
  wire  _T_1248; // @[FaultDetector.scala 334:73:@349.4]
  wire  _T_1249; // @[FaultDetector.scala 335:49:@351.4]
  wire [3:0] _T_1252; // @[FaultDetector.scala 336:50:@354.4]
  wire  _T_1254; // @[FaultDetector.scala 336:74:@355.4]
  wire [2:0] _T_1255; // @[FaultDetector.scala 337:49:@357.4]
  wire  _T_1257; // @[FaultDetector.scala 337:72:@358.4]
  wire [3:0] _T_1258; // @[FaultDetector.scala 338:48:@360.4]
  wire  _T_1260; // @[FaultDetector.scala 338:70:@361.4]
  wire [3:0] _T_1261; // @[FaultDetector.scala 340:47:@363.4]
  wire  _T_1263; // @[FaultDetector.scala 340:68:@364.4]
  wire [31:0] _T_1264; // @[FaultDetector.scala 341:49:@366.4]
  wire  _T_1266; // @[FaultDetector.scala 341:72:@367.4]
  wire [7:0] _T_1267; // @[FaultDetector.scala 342:48:@369.4]
  wire  _T_1269; // @[FaultDetector.scala 342:70:@370.4]
  wire [2:0] _T_1270; // @[FaultDetector.scala 343:49:@372.4]
  wire  _T_1272; // @[FaultDetector.scala 343:72:@373.4]
  wire [1:0] _T_1273; // @[FaultDetector.scala 344:50:@375.4]
  wire  _T_1275; // @[FaultDetector.scala 344:74:@376.4]
  wire  _T_1276; // @[FaultDetector.scala 345:49:@378.4]
  wire [3:0] _T_1279; // @[FaultDetector.scala 346:50:@381.4]
  wire  _T_1281; // @[FaultDetector.scala 346:74:@382.4]
  wire [2:0] _T_1282; // @[FaultDetector.scala 347:49:@384.4]
  wire  _T_1284; // @[FaultDetector.scala 347:72:@385.4]
  wire [3:0] _T_1285; // @[FaultDetector.scala 348:48:@387.4]
  wire  _T_1287; // @[FaultDetector.scala 348:70:@388.4]
  wire [31:0] _T_1288; // @[FaultDetector.scala 350:48:@390.4]
  wire  _T_1290; // @[FaultDetector.scala 350:70:@391.4]
  wire [3:0] _T_1291; // @[FaultDetector.scala 351:48:@393.4]
  wire  _T_1293; // @[FaultDetector.scala 351:70:@394.4]
  wire  _T_1294; // @[FaultDetector.scala 352:48:@396.4]
  wire  _T_1351; // @[FaultDetector.scala 354:46:@426.4]
  wire  _T_1352; // @[FaultDetector.scala 354:46:@427.4]
  wire  _T_1353; // @[FaultDetector.scala 354:46:@428.4]
  wire  _T_1354; // @[FaultDetector.scala 354:46:@429.4]
  wire  _T_1355; // @[FaultDetector.scala 354:46:@430.4]
  wire  _T_1356; // @[FaultDetector.scala 354:46:@431.4]
  wire  _T_1357; // @[FaultDetector.scala 354:46:@432.4]
  wire  _T_1358; // @[FaultDetector.scala 354:46:@433.4]
  wire  _T_1359; // @[FaultDetector.scala 354:46:@434.4]
  wire  _T_1360; // @[FaultDetector.scala 354:46:@435.4]
  wire  _T_1361; // @[FaultDetector.scala 354:46:@436.4]
  wire  _T_1362; // @[FaultDetector.scala 354:46:@437.4]
  wire  _T_1363; // @[FaultDetector.scala 354:46:@438.4]
  wire  _T_1364; // @[FaultDetector.scala 354:46:@439.4]
  wire  _T_1365; // @[FaultDetector.scala 354:46:@440.4]
  wire  _T_1366; // @[FaultDetector.scala 354:46:@441.4]
  wire  _T_1367; // @[FaultDetector.scala 354:46:@442.4]
  wire  _T_1368; // @[FaultDetector.scala 354:46:@443.4]
  wire  _T_1369; // @[FaultDetector.scala 354:46:@444.4]
  wire  _T_1370; // @[FaultDetector.scala 354:46:@445.4]
  wire  _T_1371; // @[FaultDetector.scala 354:46:@446.4]
  wire  _T_1372; // @[FaultDetector.scala 354:46:@447.4]
  wire  _T_1373; // @[FaultDetector.scala 354:46:@448.4]
  wire  _T_1374; // @[FaultDetector.scala 354:46:@449.4]
  wire  _T_1375; // @[FaultDetector.scala 354:46:@450.4]
  wire  _T_1376; // @[FaultDetector.scala 323:43:@452.4]
  wire  _T_1377; // @[FaultDetector.scala 324:42:@454.4]
  wire  _T_1378; // @[FaultDetector.scala 325:43:@456.4]
  wire  _T_1379; // @[FaultDetector.scala 327:42:@458.4]
  wire  _T_1380; // @[FaultDetector.scala 328:42:@460.4]
  wire [3:0] _T_1381; // @[FaultDetector.scala 330:46:@462.4]
  wire  _T_1383; // @[FaultDetector.scala 330:67:@463.4]
  wire [31:0] _T_1384; // @[FaultDetector.scala 331:48:@465.4]
  wire  _T_1386; // @[FaultDetector.scala 331:71:@466.4]
  wire [7:0] _T_1387; // @[FaultDetector.scala 332:47:@468.4]
  wire  _T_1389; // @[FaultDetector.scala 332:69:@469.4]
  wire [2:0] _T_1390; // @[FaultDetector.scala 333:48:@471.4]
  wire  _T_1392; // @[FaultDetector.scala 333:71:@472.4]
  wire [1:0] _T_1393; // @[FaultDetector.scala 334:49:@474.4]
  wire  _T_1395; // @[FaultDetector.scala 334:73:@475.4]
  wire  _T_1396; // @[FaultDetector.scala 335:49:@477.4]
  wire [3:0] _T_1399; // @[FaultDetector.scala 336:50:@480.4]
  wire  _T_1401; // @[FaultDetector.scala 336:74:@481.4]
  wire [2:0] _T_1402; // @[FaultDetector.scala 337:49:@483.4]
  wire  _T_1404; // @[FaultDetector.scala 337:72:@484.4]
  wire [3:0] _T_1405; // @[FaultDetector.scala 338:48:@486.4]
  wire  _T_1407; // @[FaultDetector.scala 338:70:@487.4]
  wire [3:0] _T_1408; // @[FaultDetector.scala 340:47:@489.4]
  wire  _T_1410; // @[FaultDetector.scala 340:68:@490.4]
  wire [31:0] _T_1411; // @[FaultDetector.scala 341:49:@492.4]
  wire  _T_1413; // @[FaultDetector.scala 341:72:@493.4]
  wire [7:0] _T_1414; // @[FaultDetector.scala 342:48:@495.4]
  wire  _T_1416; // @[FaultDetector.scala 342:70:@496.4]
  wire [2:0] _T_1417; // @[FaultDetector.scala 343:49:@498.4]
  wire  _T_1419; // @[FaultDetector.scala 343:72:@499.4]
  wire [1:0] _T_1420; // @[FaultDetector.scala 344:50:@501.4]
  wire  _T_1422; // @[FaultDetector.scala 344:74:@502.4]
  wire  _T_1423; // @[FaultDetector.scala 345:49:@504.4]
  wire [3:0] _T_1426; // @[FaultDetector.scala 346:50:@507.4]
  wire  _T_1428; // @[FaultDetector.scala 346:74:@508.4]
  wire [2:0] _T_1429; // @[FaultDetector.scala 347:49:@510.4]
  wire  _T_1431; // @[FaultDetector.scala 347:72:@511.4]
  wire [3:0] _T_1432; // @[FaultDetector.scala 348:48:@513.4]
  wire  _T_1434; // @[FaultDetector.scala 348:70:@514.4]
  wire [31:0] _T_1435; // @[FaultDetector.scala 350:48:@516.4]
  wire  _T_1437; // @[FaultDetector.scala 350:70:@517.4]
  wire [3:0] _T_1438; // @[FaultDetector.scala 351:48:@519.4]
  wire  _T_1440; // @[FaultDetector.scala 351:70:@520.4]
  wire  _T_1441; // @[FaultDetector.scala 352:48:@522.4]
  wire  _T_1498; // @[FaultDetector.scala 354:46:@552.4]
  wire  _T_1499; // @[FaultDetector.scala 354:46:@553.4]
  wire  _T_1500; // @[FaultDetector.scala 354:46:@554.4]
  wire  _T_1501; // @[FaultDetector.scala 354:46:@555.4]
  wire  _T_1502; // @[FaultDetector.scala 354:46:@556.4]
  wire  _T_1503; // @[FaultDetector.scala 354:46:@557.4]
  wire  _T_1504; // @[FaultDetector.scala 354:46:@558.4]
  wire  _T_1505; // @[FaultDetector.scala 354:46:@559.4]
  wire  _T_1506; // @[FaultDetector.scala 354:46:@560.4]
  wire  _T_1507; // @[FaultDetector.scala 354:46:@561.4]
  wire  _T_1508; // @[FaultDetector.scala 354:46:@562.4]
  wire  _T_1509; // @[FaultDetector.scala 354:46:@563.4]
  wire  _T_1510; // @[FaultDetector.scala 354:46:@564.4]
  wire  _T_1511; // @[FaultDetector.scala 354:46:@565.4]
  wire  _T_1512; // @[FaultDetector.scala 354:46:@566.4]
  wire  _T_1513; // @[FaultDetector.scala 354:46:@567.4]
  wire  _T_1514; // @[FaultDetector.scala 354:46:@568.4]
  wire  _T_1515; // @[FaultDetector.scala 354:46:@569.4]
  wire  _T_1516; // @[FaultDetector.scala 354:46:@570.4]
  wire  _T_1517; // @[FaultDetector.scala 354:46:@571.4]
  wire  _T_1518; // @[FaultDetector.scala 354:46:@572.4]
  wire  _T_1519; // @[FaultDetector.scala 354:46:@573.4]
  wire  _T_1520; // @[FaultDetector.scala 354:46:@574.4]
  wire  _T_1521; // @[FaultDetector.scala 354:46:@575.4]
  wire  _T_1522; // @[FaultDetector.scala 354:46:@576.4]
  wire  _T_1523; // @[FaultDetector.scala 323:43:@578.4]
  wire  _T_1524; // @[FaultDetector.scala 324:42:@580.4]
  wire  _T_1525; // @[FaultDetector.scala 325:43:@582.4]
  wire  _T_1526; // @[FaultDetector.scala 327:42:@584.4]
  wire  _T_1527; // @[FaultDetector.scala 328:42:@586.4]
  wire [3:0] _T_1528; // @[FaultDetector.scala 330:46:@588.4]
  wire  _T_1530; // @[FaultDetector.scala 330:67:@589.4]
  wire [31:0] _T_1531; // @[FaultDetector.scala 331:48:@591.4]
  wire  _T_1533; // @[FaultDetector.scala 331:71:@592.4]
  wire [7:0] _T_1534; // @[FaultDetector.scala 332:47:@594.4]
  wire  _T_1536; // @[FaultDetector.scala 332:69:@595.4]
  wire [2:0] _T_1537; // @[FaultDetector.scala 333:48:@597.4]
  wire  _T_1539; // @[FaultDetector.scala 333:71:@598.4]
  wire [1:0] _T_1540; // @[FaultDetector.scala 334:49:@600.4]
  wire  _T_1542; // @[FaultDetector.scala 334:73:@601.4]
  wire  _T_1543; // @[FaultDetector.scala 335:49:@603.4]
  wire [3:0] _T_1546; // @[FaultDetector.scala 336:50:@606.4]
  wire  _T_1548; // @[FaultDetector.scala 336:74:@607.4]
  wire [2:0] _T_1549; // @[FaultDetector.scala 337:49:@609.4]
  wire  _T_1551; // @[FaultDetector.scala 337:72:@610.4]
  wire [3:0] _T_1552; // @[FaultDetector.scala 338:48:@612.4]
  wire  _T_1554; // @[FaultDetector.scala 338:70:@613.4]
  wire [3:0] _T_1555; // @[FaultDetector.scala 340:47:@615.4]
  wire  _T_1557; // @[FaultDetector.scala 340:68:@616.4]
  wire [31:0] _T_1558; // @[FaultDetector.scala 341:49:@618.4]
  wire  _T_1560; // @[FaultDetector.scala 341:72:@619.4]
  wire [7:0] _T_1561; // @[FaultDetector.scala 342:48:@621.4]
  wire  _T_1563; // @[FaultDetector.scala 342:70:@622.4]
  wire [2:0] _T_1564; // @[FaultDetector.scala 343:49:@624.4]
  wire  _T_1566; // @[FaultDetector.scala 343:72:@625.4]
  wire [1:0] _T_1567; // @[FaultDetector.scala 344:50:@627.4]
  wire  _T_1569; // @[FaultDetector.scala 344:74:@628.4]
  wire  _T_1570; // @[FaultDetector.scala 345:49:@630.4]
  wire [3:0] _T_1573; // @[FaultDetector.scala 346:50:@633.4]
  wire  _T_1575; // @[FaultDetector.scala 346:74:@634.4]
  wire [2:0] _T_1576; // @[FaultDetector.scala 347:49:@636.4]
  wire  _T_1578; // @[FaultDetector.scala 347:72:@637.4]
  wire [3:0] _T_1579; // @[FaultDetector.scala 348:48:@639.4]
  wire  _T_1581; // @[FaultDetector.scala 348:70:@640.4]
  wire [31:0] _T_1582; // @[FaultDetector.scala 350:48:@642.4]
  wire  _T_1584; // @[FaultDetector.scala 350:70:@643.4]
  wire [3:0] _T_1585; // @[FaultDetector.scala 351:48:@645.4]
  wire  _T_1587; // @[FaultDetector.scala 351:70:@646.4]
  wire  _T_1588; // @[FaultDetector.scala 352:48:@648.4]
  wire  _T_1645; // @[FaultDetector.scala 354:46:@678.4]
  wire  _T_1646; // @[FaultDetector.scala 354:46:@679.4]
  wire  _T_1647; // @[FaultDetector.scala 354:46:@680.4]
  wire  _T_1648; // @[FaultDetector.scala 354:46:@681.4]
  wire  _T_1649; // @[FaultDetector.scala 354:46:@682.4]
  wire  _T_1650; // @[FaultDetector.scala 354:46:@683.4]
  wire  _T_1651; // @[FaultDetector.scala 354:46:@684.4]
  wire  _T_1652; // @[FaultDetector.scala 354:46:@685.4]
  wire  _T_1653; // @[FaultDetector.scala 354:46:@686.4]
  wire  _T_1654; // @[FaultDetector.scala 354:46:@687.4]
  wire  _T_1655; // @[FaultDetector.scala 354:46:@688.4]
  wire  _T_1656; // @[FaultDetector.scala 354:46:@689.4]
  wire  _T_1657; // @[FaultDetector.scala 354:46:@690.4]
  wire  _T_1658; // @[FaultDetector.scala 354:46:@691.4]
  wire  _T_1659; // @[FaultDetector.scala 354:46:@692.4]
  wire  _T_1660; // @[FaultDetector.scala 354:46:@693.4]
  wire  _T_1661; // @[FaultDetector.scala 354:46:@694.4]
  wire  _T_1662; // @[FaultDetector.scala 354:46:@695.4]
  wire  _T_1663; // @[FaultDetector.scala 354:46:@696.4]
  wire  _T_1664; // @[FaultDetector.scala 354:46:@697.4]
  wire  _T_1665; // @[FaultDetector.scala 354:46:@698.4]
  wire  _T_1666; // @[FaultDetector.scala 354:46:@699.4]
  wire  _T_1667; // @[FaultDetector.scala 354:46:@700.4]
  wire  _T_1668; // @[FaultDetector.scala 354:46:@701.4]
  wire  _T_1669; // @[FaultDetector.scala 354:46:@702.4]
  wire [1:0] _T_1672; // @[Cat.scala 30:58:@704.4]
  wire [2:0] _T_1673; // @[Cat.scala 30:58:@705.4]
  wire [3:0] _T_1674; // @[Cat.scala 30:58:@706.4]
  wire [3:0] invalid; // @[FaultDetector.scala 358:8:@707.4]
  reg [2:0] invalid_reg; // @[FaultDetector.scala 426:28:@708.4]
  reg [31:0] _RAND_223;
  reg [2:0] faulty_cpu; // @[FaultDetector.scala 427:27:@709.4]
  reg [31:0] _RAND_224;
  reg  reset_logic_reg; // @[FaultDetector.scala 429:32:@710.4]
  reg [31:0] _RAND_225;
  reg  cpu_back_online_reg; // @[FaultDetector.scala 431:36:@711.4]
  reg [31:0] _RAND_226;
  wire  ack_back_online; // @[FaultDetector.scala 432:29:@712.4]
  wire  _GEN_0; // @[FaultDetector.scala 434:28:@714.4]
  wire [2:0] _GEN_5; // @[FaultDetector.scala 434:28:@714.4]
  wire  _T_1693; // @[FaultDetector.scala 444:18:@724.6]
  wire  _GEN_7; // @[FaultDetector.scala 444:27:@725.6]
  wire  _GEN_8; // @[FaultDetector.scala 444:27:@725.6]
  wire  _GEN_9; // @[FaultDetector.scala 443:25:@723.4]
  wire  _GEN_10; // @[FaultDetector.scala 443:25:@723.4]
  wire  _GEN_11; // @[FaultDetector.scala 450:25:@730.4]
  wire  _T_1698; // @[FaultDetector.scala 456:16:@734.4]
  wire  _T_1701; // @[FaultDetector.scala 456:27:@736.4]
  wire  _T_1702; // @[FaultDetector.scala 456:24:@737.4]
  wire [3:0] _GEN_12; // @[FaultDetector.scala 456:52:@738.4]
  wire  _T_1704; // @[FaultDetector.scala 460:20:@741.4]
  wire [2:0] _T_1705; // @[FaultDetector.scala 462:21:@743.6]
  wire [2:0] _GEN_13; // @[FaultDetector.scala 460:29:@742.4]
  wire  _T_1709; // @[FaultDetector.scala 473:30:@753.4]
  wire  _T_1710; // @[FaultDetector.scala 473:30:@757.4]
  wire  _T_1711; // @[FaultDetector.scala 473:30:@761.4]
  wire  invalid_bool_0; // @[FaultDetector.scala 477:33:@764.4]
  wire  invalid_bool_1; // @[FaultDetector.scala 477:33:@765.4]
  wire  invalid_bool_2; // @[FaultDetector.scala 477:33:@766.4]
  wire  _T_1713; // @[FaultDetector.scala 121:8:@767.4]
  wire  _GEN_15; // @[FaultDetector.scala 125:21:@772.6]
  wire  _GEN_16; // @[FaultDetector.scala 125:21:@772.6]
  wire  _GEN_17; // @[FaultDetector.scala 125:21:@772.6]
  wire  _GEN_18; // @[FaultDetector.scala 125:21:@772.6]
  wire [3:0] _GEN_19; // @[FaultDetector.scala 125:21:@772.6]
  wire [1:0] _GEN_20; // @[FaultDetector.scala 125:21:@772.6]
  wire  _GEN_21; // @[FaultDetector.scala 125:21:@772.6]
  wire [3:0] _GEN_22; // @[FaultDetector.scala 125:21:@772.6]
  wire [1:0] _GEN_23; // @[FaultDetector.scala 125:21:@772.6]
  wire  _GEN_24; // @[FaultDetector.scala 125:21:@772.6]
  wire [31:0] _GEN_25; // @[FaultDetector.scala 125:21:@772.6]
  wire  _GEN_26; // @[FaultDetector.scala 121:15:@768.4]
  wire  _GEN_37; // @[FaultDetector.scala 121:15:@768.4]
  wire  _GEN_43; // @[FaultDetector.scala 121:15:@768.4]
  wire [3:0] _GEN_44; // @[FaultDetector.scala 121:15:@768.4]
  wire [1:0] _GEN_45; // @[FaultDetector.scala 121:15:@768.4]
  wire  _GEN_46; // @[FaultDetector.scala 121:15:@768.4]
  wire  _GEN_58; // @[FaultDetector.scala 121:15:@768.4]
  wire [3:0] _GEN_59; // @[FaultDetector.scala 121:15:@768.4]
  wire [31:0] _GEN_60; // @[FaultDetector.scala 121:15:@768.4]
  wire [1:0] _GEN_61; // @[FaultDetector.scala 121:15:@768.4]
  wire  _GEN_62; // @[FaultDetector.scala 121:15:@768.4]
  wire  _GEN_63; // @[FaultDetector.scala 121:15:@768.4]
  wire  _GEN_64; // @[FaultDetector.scala 121:15:@768.4]
  wire [3:0] _GEN_65; // @[FaultDetector.scala 121:15:@768.4]
  wire [31:0] _GEN_66; // @[FaultDetector.scala 121:15:@768.4]
  wire [7:0] _GEN_67; // @[FaultDetector.scala 121:15:@768.4]
  wire [2:0] _GEN_68; // @[FaultDetector.scala 121:15:@768.4]
  wire [1:0] _GEN_69; // @[FaultDetector.scala 121:15:@768.4]
  wire  _GEN_70; // @[FaultDetector.scala 121:15:@768.4]
  wire [3:0] _GEN_71; // @[FaultDetector.scala 121:15:@768.4]
  wire [2:0] _GEN_72; // @[FaultDetector.scala 121:15:@768.4]
  wire [3:0] _GEN_73; // @[FaultDetector.scala 121:15:@768.4]
  wire  _GEN_74; // @[FaultDetector.scala 121:15:@768.4]
  wire  _GEN_75; // @[FaultDetector.scala 121:15:@768.4]
  wire [31:0] _GEN_76; // @[FaultDetector.scala 121:15:@768.4]
  wire [3:0] _GEN_77; // @[FaultDetector.scala 121:15:@768.4]
  wire  _GEN_78; // @[FaultDetector.scala 121:15:@768.4]
  wire  _GEN_79; // @[FaultDetector.scala 121:15:@768.4]
  wire  _GEN_80; // @[FaultDetector.scala 121:15:@768.4]
  wire [3:0] _GEN_81; // @[FaultDetector.scala 121:15:@768.4]
  wire [1:0] _GEN_82; // @[FaultDetector.scala 121:15:@768.4]
  wire  _GEN_83; // @[FaultDetector.scala 121:15:@768.4]
  wire  _GEN_84; // @[FaultDetector.scala 121:15:@768.4]
  wire [3:0] _GEN_85; // @[FaultDetector.scala 121:15:@768.4]
  wire [31:0] _GEN_86; // @[FaultDetector.scala 121:15:@768.4]
  wire [7:0] _GEN_87; // @[FaultDetector.scala 121:15:@768.4]
  wire [2:0] _GEN_88; // @[FaultDetector.scala 121:15:@768.4]
  wire [1:0] _GEN_89; // @[FaultDetector.scala 121:15:@768.4]
  wire  _GEN_90; // @[FaultDetector.scala 121:15:@768.4]
  wire [3:0] _GEN_91; // @[FaultDetector.scala 121:15:@768.4]
  wire [2:0] _GEN_92; // @[FaultDetector.scala 121:15:@768.4]
  wire [3:0] _GEN_93; // @[FaultDetector.scala 121:15:@768.4]
  wire  _GEN_94; // @[FaultDetector.scala 121:15:@768.4]
  wire  _GEN_95; // @[FaultDetector.scala 121:15:@768.4]
  wire [3:0] _GEN_96; // @[FaultDetector.scala 121:15:@768.4]
  wire [31:0] _GEN_97; // @[FaultDetector.scala 121:15:@768.4]
  wire [1:0] _GEN_98; // @[FaultDetector.scala 121:15:@768.4]
  wire  _GEN_99; // @[FaultDetector.scala 121:15:@768.4]
  wire  _T_1726; // @[FaultDetector.scala 121:8:@790.4]
  wire  _GEN_137; // @[FaultDetector.scala 125:21:@795.6]
  wire  _GEN_138; // @[FaultDetector.scala 125:21:@795.6]
  wire  _GEN_139; // @[FaultDetector.scala 125:21:@795.6]
  wire  _GEN_140; // @[FaultDetector.scala 125:21:@795.6]
  wire [3:0] _GEN_141; // @[FaultDetector.scala 125:21:@795.6]
  wire [1:0] _GEN_142; // @[FaultDetector.scala 125:21:@795.6]
  wire  _GEN_143; // @[FaultDetector.scala 125:21:@795.6]
  wire [3:0] _GEN_144; // @[FaultDetector.scala 125:21:@795.6]
  wire [1:0] _GEN_145; // @[FaultDetector.scala 125:21:@795.6]
  wire  _GEN_146; // @[FaultDetector.scala 125:21:@795.6]
  wire [31:0] _GEN_147; // @[FaultDetector.scala 125:21:@795.6]
  wire  _GEN_148; // @[FaultDetector.scala 121:15:@791.4]
  wire  _GEN_159; // @[FaultDetector.scala 121:15:@791.4]
  wire  _GEN_165; // @[FaultDetector.scala 121:15:@791.4]
  wire [3:0] _GEN_166; // @[FaultDetector.scala 121:15:@791.4]
  wire [1:0] _GEN_167; // @[FaultDetector.scala 121:15:@791.4]
  wire  _GEN_168; // @[FaultDetector.scala 121:15:@791.4]
  wire  _GEN_180; // @[FaultDetector.scala 121:15:@791.4]
  wire [3:0] _GEN_181; // @[FaultDetector.scala 121:15:@791.4]
  wire [31:0] _GEN_182; // @[FaultDetector.scala 121:15:@791.4]
  wire [1:0] _GEN_183; // @[FaultDetector.scala 121:15:@791.4]
  wire  _GEN_184; // @[FaultDetector.scala 121:15:@791.4]
  wire  _GEN_185; // @[FaultDetector.scala 121:15:@791.4]
  wire  _GEN_186; // @[FaultDetector.scala 121:15:@791.4]
  wire [3:0] _GEN_187; // @[FaultDetector.scala 121:15:@791.4]
  wire [31:0] _GEN_188; // @[FaultDetector.scala 121:15:@791.4]
  wire [7:0] _GEN_189; // @[FaultDetector.scala 121:15:@791.4]
  wire [2:0] _GEN_190; // @[FaultDetector.scala 121:15:@791.4]
  wire [1:0] _GEN_191; // @[FaultDetector.scala 121:15:@791.4]
  wire  _GEN_192; // @[FaultDetector.scala 121:15:@791.4]
  wire [3:0] _GEN_193; // @[FaultDetector.scala 121:15:@791.4]
  wire [2:0] _GEN_194; // @[FaultDetector.scala 121:15:@791.4]
  wire [3:0] _GEN_195; // @[FaultDetector.scala 121:15:@791.4]
  wire  _GEN_196; // @[FaultDetector.scala 121:15:@791.4]
  wire  _GEN_197; // @[FaultDetector.scala 121:15:@791.4]
  wire [31:0] _GEN_198; // @[FaultDetector.scala 121:15:@791.4]
  wire [3:0] _GEN_199; // @[FaultDetector.scala 121:15:@791.4]
  wire  _GEN_200; // @[FaultDetector.scala 121:15:@791.4]
  wire  _GEN_201; // @[FaultDetector.scala 121:15:@791.4]
  wire  _GEN_202; // @[FaultDetector.scala 121:15:@791.4]
  wire [3:0] _GEN_203; // @[FaultDetector.scala 121:15:@791.4]
  wire [1:0] _GEN_204; // @[FaultDetector.scala 121:15:@791.4]
  wire  _GEN_205; // @[FaultDetector.scala 121:15:@791.4]
  wire  _GEN_206; // @[FaultDetector.scala 121:15:@791.4]
  wire [3:0] _GEN_207; // @[FaultDetector.scala 121:15:@791.4]
  wire [31:0] _GEN_208; // @[FaultDetector.scala 121:15:@791.4]
  wire [7:0] _GEN_209; // @[FaultDetector.scala 121:15:@791.4]
  wire [2:0] _GEN_210; // @[FaultDetector.scala 121:15:@791.4]
  wire [1:0] _GEN_211; // @[FaultDetector.scala 121:15:@791.4]
  wire  _GEN_212; // @[FaultDetector.scala 121:15:@791.4]
  wire [3:0] _GEN_213; // @[FaultDetector.scala 121:15:@791.4]
  wire [2:0] _GEN_214; // @[FaultDetector.scala 121:15:@791.4]
  wire [3:0] _GEN_215; // @[FaultDetector.scala 121:15:@791.4]
  wire  _GEN_216; // @[FaultDetector.scala 121:15:@791.4]
  wire  _GEN_217; // @[FaultDetector.scala 121:15:@791.4]
  wire [3:0] _GEN_218; // @[FaultDetector.scala 121:15:@791.4]
  wire [31:0] _GEN_219; // @[FaultDetector.scala 121:15:@791.4]
  wire [1:0] _GEN_220; // @[FaultDetector.scala 121:15:@791.4]
  wire  _GEN_221; // @[FaultDetector.scala 121:15:@791.4]
  wire  _T_1739; // @[FaultDetector.scala 121:8:@813.4]
  wire  _GEN_259; // @[FaultDetector.scala 125:21:@818.6]
  wire  _GEN_260; // @[FaultDetector.scala 125:21:@818.6]
  wire  _GEN_261; // @[FaultDetector.scala 125:21:@818.6]
  wire  _GEN_262; // @[FaultDetector.scala 125:21:@818.6]
  wire [3:0] _GEN_263; // @[FaultDetector.scala 125:21:@818.6]
  wire [1:0] _GEN_264; // @[FaultDetector.scala 125:21:@818.6]
  wire  _GEN_265; // @[FaultDetector.scala 125:21:@818.6]
  wire [3:0] _GEN_266; // @[FaultDetector.scala 125:21:@818.6]
  wire [1:0] _GEN_267; // @[FaultDetector.scala 125:21:@818.6]
  wire  _GEN_268; // @[FaultDetector.scala 125:21:@818.6]
  wire [31:0] _GEN_269; // @[FaultDetector.scala 125:21:@818.6]
  wire  _GEN_270; // @[FaultDetector.scala 121:15:@814.4]
  wire  _GEN_281; // @[FaultDetector.scala 121:15:@814.4]
  wire  _GEN_287; // @[FaultDetector.scala 121:15:@814.4]
  wire [3:0] _GEN_288; // @[FaultDetector.scala 121:15:@814.4]
  wire [1:0] _GEN_289; // @[FaultDetector.scala 121:15:@814.4]
  wire  _GEN_290; // @[FaultDetector.scala 121:15:@814.4]
  wire  _GEN_302; // @[FaultDetector.scala 121:15:@814.4]
  wire [3:0] _GEN_303; // @[FaultDetector.scala 121:15:@814.4]
  wire [31:0] _GEN_304; // @[FaultDetector.scala 121:15:@814.4]
  wire [1:0] _GEN_305; // @[FaultDetector.scala 121:15:@814.4]
  wire  _GEN_306; // @[FaultDetector.scala 121:15:@814.4]
  wire  _GEN_307; // @[FaultDetector.scala 121:15:@814.4]
  wire  _GEN_308; // @[FaultDetector.scala 121:15:@814.4]
  wire [3:0] _GEN_309; // @[FaultDetector.scala 121:15:@814.4]
  wire [31:0] _GEN_310; // @[FaultDetector.scala 121:15:@814.4]
  wire [7:0] _GEN_311; // @[FaultDetector.scala 121:15:@814.4]
  wire [2:0] _GEN_312; // @[FaultDetector.scala 121:15:@814.4]
  wire [1:0] _GEN_313; // @[FaultDetector.scala 121:15:@814.4]
  wire  _GEN_314; // @[FaultDetector.scala 121:15:@814.4]
  wire [3:0] _GEN_315; // @[FaultDetector.scala 121:15:@814.4]
  wire [2:0] _GEN_316; // @[FaultDetector.scala 121:15:@814.4]
  wire [3:0] _GEN_317; // @[FaultDetector.scala 121:15:@814.4]
  wire  _GEN_318; // @[FaultDetector.scala 121:15:@814.4]
  wire  _GEN_319; // @[FaultDetector.scala 121:15:@814.4]
  wire [31:0] _GEN_320; // @[FaultDetector.scala 121:15:@814.4]
  wire [3:0] _GEN_321; // @[FaultDetector.scala 121:15:@814.4]
  wire  _GEN_322; // @[FaultDetector.scala 121:15:@814.4]
  wire  _GEN_323; // @[FaultDetector.scala 121:15:@814.4]
  wire  _GEN_324; // @[FaultDetector.scala 121:15:@814.4]
  wire [3:0] _GEN_325; // @[FaultDetector.scala 121:15:@814.4]
  wire [1:0] _GEN_326; // @[FaultDetector.scala 121:15:@814.4]
  wire  _GEN_327; // @[FaultDetector.scala 121:15:@814.4]
  wire  _GEN_328; // @[FaultDetector.scala 121:15:@814.4]
  wire [3:0] _GEN_329; // @[FaultDetector.scala 121:15:@814.4]
  wire [31:0] _GEN_330; // @[FaultDetector.scala 121:15:@814.4]
  wire [7:0] _GEN_331; // @[FaultDetector.scala 121:15:@814.4]
  wire [2:0] _GEN_332; // @[FaultDetector.scala 121:15:@814.4]
  wire [1:0] _GEN_333; // @[FaultDetector.scala 121:15:@814.4]
  wire  _GEN_334; // @[FaultDetector.scala 121:15:@814.4]
  wire [3:0] _GEN_335; // @[FaultDetector.scala 121:15:@814.4]
  wire [2:0] _GEN_336; // @[FaultDetector.scala 121:15:@814.4]
  wire [3:0] _GEN_337; // @[FaultDetector.scala 121:15:@814.4]
  wire  _GEN_338; // @[FaultDetector.scala 121:15:@814.4]
  wire  _GEN_339; // @[FaultDetector.scala 121:15:@814.4]
  wire [3:0] _GEN_340; // @[FaultDetector.scala 121:15:@814.4]
  wire [31:0] _GEN_341; // @[FaultDetector.scala 121:15:@814.4]
  wire [1:0] _GEN_342; // @[FaultDetector.scala 121:15:@814.4]
  wire  _GEN_343; // @[FaultDetector.scala 121:15:@814.4]
  wire  _T_1752; // @[FaultDetector.scala 177:24:@869.4]
  wire  _T_1753; // @[FaultDetector.scala 179:56:@871.6]
  wire  _T_1754; // @[FaultDetector.scala 180:56:@873.6]
  wire  _T_1755; // @[FaultDetector.scala 181:56:@875.6]
  wire  _T_1756; // @[FaultDetector.scala 183:54:@877.6]
  wire  _T_1757; // @[FaultDetector.scala 184:54:@879.6]
  wire [3:0] _T_1758; // @[FaultDetector.scala 186:66:@881.6]
  wire [31:0] _T_1759; // @[FaultDetector.scala 187:66:@883.6]
  wire [7:0] _T_1760; // @[FaultDetector.scala 188:66:@885.6]
  wire [2:0] _T_1761; // @[FaultDetector.scala 189:66:@887.6]
  wire [1:0] _T_1762; // @[FaultDetector.scala 190:66:@889.6]
  wire  _T_1763; // @[FaultDetector.scala 191:66:@891.6]
  wire [3:0] _T_1764; // @[FaultDetector.scala 192:66:@893.6]
  wire [2:0] _T_1765; // @[FaultDetector.scala 193:66:@895.6]
  wire [3:0] _T_1766; // @[FaultDetector.scala 194:66:@897.6]
  wire [3:0] _T_1767; // @[FaultDetector.scala 196:66:@899.6]
  wire [31:0] _T_1768; // @[FaultDetector.scala 197:66:@901.6]
  wire [7:0] _T_1769; // @[FaultDetector.scala 198:66:@903.6]
  wire [2:0] _T_1770; // @[FaultDetector.scala 199:66:@905.6]
  wire [1:0] _T_1771; // @[FaultDetector.scala 200:66:@907.6]
  wire  _T_1772; // @[FaultDetector.scala 201:66:@909.6]
  wire [3:0] _T_1773; // @[FaultDetector.scala 202:66:@911.6]
  wire [2:0] _T_1774; // @[FaultDetector.scala 203:66:@913.6]
  wire [3:0] _T_1775; // @[FaultDetector.scala 204:66:@915.6]
  wire [31:0] _T_1776; // @[FaultDetector.scala 206:62:@917.6]
  wire [3:0] _T_1777; // @[FaultDetector.scala 207:62:@919.6]
  wire  _T_1778; // @[FaultDetector.scala 208:62:@921.6]
  wire  _T_1780; // @[FaultDetector.scala 210:30:@925.6]
  wire  _T_1781; // @[FaultDetector.scala 212:56:@927.8]
  wire  _T_1782; // @[FaultDetector.scala 213:56:@929.8]
  wire  _T_1783; // @[FaultDetector.scala 214:56:@931.8]
  wire  _T_1784; // @[FaultDetector.scala 216:54:@933.8]
  wire  _T_1785; // @[FaultDetector.scala 217:54:@935.8]
  wire [3:0] _T_1786; // @[FaultDetector.scala 219:66:@937.8]
  wire [31:0] _T_1787; // @[FaultDetector.scala 220:66:@939.8]
  wire [7:0] _T_1788; // @[FaultDetector.scala 221:66:@941.8]
  wire [2:0] _T_1789; // @[FaultDetector.scala 222:66:@943.8]
  wire [1:0] _T_1790; // @[FaultDetector.scala 223:66:@945.8]
  wire  _T_1791; // @[FaultDetector.scala 224:66:@947.8]
  wire [3:0] _T_1792; // @[FaultDetector.scala 225:66:@949.8]
  wire [2:0] _T_1793; // @[FaultDetector.scala 226:66:@951.8]
  wire [3:0] _T_1794; // @[FaultDetector.scala 227:66:@953.8]
  wire [3:0] _T_1795; // @[FaultDetector.scala 229:66:@955.8]
  wire [31:0] _T_1796; // @[FaultDetector.scala 230:66:@957.8]
  wire [7:0] _T_1797; // @[FaultDetector.scala 231:66:@959.8]
  wire [2:0] _T_1798; // @[FaultDetector.scala 232:66:@961.8]
  wire [1:0] _T_1799; // @[FaultDetector.scala 233:66:@963.8]
  wire  _T_1800; // @[FaultDetector.scala 234:66:@965.8]
  wire [3:0] _T_1801; // @[FaultDetector.scala 235:66:@967.8]
  wire [2:0] _T_1802; // @[FaultDetector.scala 236:66:@969.8]
  wire [3:0] _T_1803; // @[FaultDetector.scala 237:66:@971.8]
  wire [31:0] _T_1804; // @[FaultDetector.scala 239:62:@973.8]
  wire [3:0] _T_1805; // @[FaultDetector.scala 240:62:@975.8]
  wire  _T_1806; // @[FaultDetector.scala 241:62:@977.8]
  wire  _T_1808; // @[FaultDetector.scala 243:30:@981.8]
  wire  _T_1809; // @[FaultDetector.scala 245:56:@983.10]
  wire  _T_1810; // @[FaultDetector.scala 246:56:@985.10]
  wire  _T_1811; // @[FaultDetector.scala 247:56:@987.10]
  wire  _T_1812; // @[FaultDetector.scala 249:54:@989.10]
  wire  _T_1813; // @[FaultDetector.scala 250:54:@991.10]
  wire [3:0] _T_1814; // @[FaultDetector.scala 252:66:@993.10]
  wire [31:0] _T_1815; // @[FaultDetector.scala 253:66:@995.10]
  wire [7:0] _T_1816; // @[FaultDetector.scala 254:66:@997.10]
  wire [2:0] _T_1817; // @[FaultDetector.scala 255:66:@999.10]
  wire [1:0] _T_1818; // @[FaultDetector.scala 256:66:@1001.10]
  wire  _T_1819; // @[FaultDetector.scala 257:66:@1003.10]
  wire [3:0] _T_1820; // @[FaultDetector.scala 258:66:@1005.10]
  wire [2:0] _T_1821; // @[FaultDetector.scala 259:66:@1007.10]
  wire [3:0] _T_1822; // @[FaultDetector.scala 260:66:@1009.10]
  wire [3:0] _T_1823; // @[FaultDetector.scala 262:66:@1011.10]
  wire [31:0] _T_1824; // @[FaultDetector.scala 263:66:@1013.10]
  wire [7:0] _T_1825; // @[FaultDetector.scala 264:66:@1015.10]
  wire [2:0] _T_1826; // @[FaultDetector.scala 265:66:@1017.10]
  wire [1:0] _T_1827; // @[FaultDetector.scala 266:66:@1019.10]
  wire  _T_1828; // @[FaultDetector.scala 267:66:@1021.10]
  wire [3:0] _T_1829; // @[FaultDetector.scala 268:66:@1023.10]
  wire [2:0] _T_1830; // @[FaultDetector.scala 269:66:@1025.10]
  wire [3:0] _T_1831; // @[FaultDetector.scala 270:66:@1027.10]
  wire [31:0] _T_1832; // @[FaultDetector.scala 272:62:@1029.10]
  wire [3:0] _T_1833; // @[FaultDetector.scala 273:62:@1031.10]
  wire  _T_1834; // @[FaultDetector.scala 274:62:@1033.10]
  wire  _T_1838; // @[FaultDetector.scala 279:80:@1039.10]
  wire  _T_1842; // @[FaultDetector.scala 280:80:@1043.10]
  wire  _T_1846; // @[FaultDetector.scala 281:80:@1047.10]
  wire  _T_1850; // @[FaultDetector.scala 283:79:@1051.10]
  wire  _T_1854; // @[FaultDetector.scala 284:79:@1055.10]
  wire [3:0] _T_1858; // @[FaultDetector.scala 286:81:@1059.10]
  wire [31:0] _T_1862; // @[FaultDetector.scala 287:81:@1063.10]
  wire [7:0] _T_1866; // @[FaultDetector.scala 288:81:@1067.10]
  wire [2:0] _T_1870; // @[FaultDetector.scala 289:81:@1071.10]
  wire [1:0] _T_1874; // @[FaultDetector.scala 290:81:@1075.10]
  wire  _T_1878; // @[FaultDetector.scala 291:81:@1079.10]
  wire [3:0] _T_1882; // @[FaultDetector.scala 292:81:@1083.10]
  wire [2:0] _T_1886; // @[FaultDetector.scala 293:81:@1087.10]
  wire [3:0] _T_1890; // @[FaultDetector.scala 294:81:@1091.10]
  wire [3:0] _T_1894; // @[FaultDetector.scala 296:81:@1095.10]
  wire [31:0] _T_1898; // @[FaultDetector.scala 297:81:@1099.10]
  wire [7:0] _T_1902; // @[FaultDetector.scala 298:81:@1103.10]
  wire [2:0] _T_1906; // @[FaultDetector.scala 299:81:@1107.10]
  wire [1:0] _T_1910; // @[FaultDetector.scala 300:81:@1111.10]
  wire  _T_1914; // @[FaultDetector.scala 301:81:@1115.10]
  wire [3:0] _T_1918; // @[FaultDetector.scala 302:81:@1119.10]
  wire [2:0] _T_1922; // @[FaultDetector.scala 303:81:@1123.10]
  wire [3:0] _T_1926; // @[FaultDetector.scala 304:81:@1127.10]
  wire [31:0] _T_1930; // @[FaultDetector.scala 306:79:@1131.10]
  wire [3:0] _T_1934; // @[FaultDetector.scala 307:79:@1135.10]
  wire  _T_1938; // @[FaultDetector.scala 308:79:@1139.10]
  wire  _GEN_381; // @[FaultDetector.scala 243:40:@982.8]
  wire  _GEN_382; // @[FaultDetector.scala 243:40:@982.8]
  wire  _GEN_383; // @[FaultDetector.scala 243:40:@982.8]
  wire  _GEN_384; // @[FaultDetector.scala 243:40:@982.8]
  wire  _GEN_385; // @[FaultDetector.scala 243:40:@982.8]
  wire [3:0] _GEN_386; // @[FaultDetector.scala 243:40:@982.8]
  wire [31:0] _GEN_387; // @[FaultDetector.scala 243:40:@982.8]
  wire [7:0] _GEN_388; // @[FaultDetector.scala 243:40:@982.8]
  wire [2:0] _GEN_389; // @[FaultDetector.scala 243:40:@982.8]
  wire [1:0] _GEN_390; // @[FaultDetector.scala 243:40:@982.8]
  wire  _GEN_391; // @[FaultDetector.scala 243:40:@982.8]
  wire [3:0] _GEN_392; // @[FaultDetector.scala 243:40:@982.8]
  wire [2:0] _GEN_393; // @[FaultDetector.scala 243:40:@982.8]
  wire [3:0] _GEN_394; // @[FaultDetector.scala 243:40:@982.8]
  wire [3:0] _GEN_395; // @[FaultDetector.scala 243:40:@982.8]
  wire [31:0] _GEN_396; // @[FaultDetector.scala 243:40:@982.8]
  wire [7:0] _GEN_397; // @[FaultDetector.scala 243:40:@982.8]
  wire [2:0] _GEN_398; // @[FaultDetector.scala 243:40:@982.8]
  wire [1:0] _GEN_399; // @[FaultDetector.scala 243:40:@982.8]
  wire  _GEN_400; // @[FaultDetector.scala 243:40:@982.8]
  wire [3:0] _GEN_401; // @[FaultDetector.scala 243:40:@982.8]
  wire [2:0] _GEN_402; // @[FaultDetector.scala 243:40:@982.8]
  wire [3:0] _GEN_403; // @[FaultDetector.scala 243:40:@982.8]
  wire [31:0] _GEN_404; // @[FaultDetector.scala 243:40:@982.8]
  wire [3:0] _GEN_405; // @[FaultDetector.scala 243:40:@982.8]
  wire  _GEN_406; // @[FaultDetector.scala 243:40:@982.8]
  wire  _GEN_407; // @[FaultDetector.scala 210:40:@926.6]
  wire  _GEN_408; // @[FaultDetector.scala 210:40:@926.6]
  wire  _GEN_409; // @[FaultDetector.scala 210:40:@926.6]
  wire  _GEN_410; // @[FaultDetector.scala 210:40:@926.6]
  wire  _GEN_411; // @[FaultDetector.scala 210:40:@926.6]
  wire [3:0] _GEN_412; // @[FaultDetector.scala 210:40:@926.6]
  wire [31:0] _GEN_413; // @[FaultDetector.scala 210:40:@926.6]
  wire [7:0] _GEN_414; // @[FaultDetector.scala 210:40:@926.6]
  wire [2:0] _GEN_415; // @[FaultDetector.scala 210:40:@926.6]
  wire [1:0] _GEN_416; // @[FaultDetector.scala 210:40:@926.6]
  wire  _GEN_417; // @[FaultDetector.scala 210:40:@926.6]
  wire [3:0] _GEN_418; // @[FaultDetector.scala 210:40:@926.6]
  wire [2:0] _GEN_419; // @[FaultDetector.scala 210:40:@926.6]
  wire [3:0] _GEN_420; // @[FaultDetector.scala 210:40:@926.6]
  wire [3:0] _GEN_421; // @[FaultDetector.scala 210:40:@926.6]
  wire [31:0] _GEN_422; // @[FaultDetector.scala 210:40:@926.6]
  wire [7:0] _GEN_423; // @[FaultDetector.scala 210:40:@926.6]
  wire [2:0] _GEN_424; // @[FaultDetector.scala 210:40:@926.6]
  wire [1:0] _GEN_425; // @[FaultDetector.scala 210:40:@926.6]
  wire  _GEN_426; // @[FaultDetector.scala 210:40:@926.6]
  wire [3:0] _GEN_427; // @[FaultDetector.scala 210:40:@926.6]
  wire [2:0] _GEN_428; // @[FaultDetector.scala 210:40:@926.6]
  wire [3:0] _GEN_429; // @[FaultDetector.scala 210:40:@926.6]
  wire [31:0] _GEN_430; // @[FaultDetector.scala 210:40:@926.6]
  wire [3:0] _GEN_431; // @[FaultDetector.scala 210:40:@926.6]
  wire  _GEN_432; // @[FaultDetector.scala 210:40:@926.6]
  wire  _GEN_433; // @[FaultDetector.scala 177:34:@870.4]
  wire  _GEN_434; // @[FaultDetector.scala 177:34:@870.4]
  wire  _GEN_435; // @[FaultDetector.scala 177:34:@870.4]
  wire  _GEN_436; // @[FaultDetector.scala 177:34:@870.4]
  wire  _GEN_437; // @[FaultDetector.scala 177:34:@870.4]
  wire [3:0] _GEN_438; // @[FaultDetector.scala 177:34:@870.4]
  wire [31:0] _GEN_439; // @[FaultDetector.scala 177:34:@870.4]
  wire [7:0] _GEN_440; // @[FaultDetector.scala 177:34:@870.4]
  wire [2:0] _GEN_441; // @[FaultDetector.scala 177:34:@870.4]
  wire [1:0] _GEN_442; // @[FaultDetector.scala 177:34:@870.4]
  wire  _GEN_443; // @[FaultDetector.scala 177:34:@870.4]
  wire [3:0] _GEN_444; // @[FaultDetector.scala 177:34:@870.4]
  wire [2:0] _GEN_445; // @[FaultDetector.scala 177:34:@870.4]
  wire [3:0] _GEN_446; // @[FaultDetector.scala 177:34:@870.4]
  wire [3:0] _GEN_447; // @[FaultDetector.scala 177:34:@870.4]
  wire [31:0] _GEN_448; // @[FaultDetector.scala 177:34:@870.4]
  wire [7:0] _GEN_449; // @[FaultDetector.scala 177:34:@870.4]
  wire [2:0] _GEN_450; // @[FaultDetector.scala 177:34:@870.4]
  wire [1:0] _GEN_451; // @[FaultDetector.scala 177:34:@870.4]
  wire  _GEN_452; // @[FaultDetector.scala 177:34:@870.4]
  wire [3:0] _GEN_453; // @[FaultDetector.scala 177:34:@870.4]
  wire [2:0] _GEN_454; // @[FaultDetector.scala 177:34:@870.4]
  wire [3:0] _GEN_455; // @[FaultDetector.scala 177:34:@870.4]
  wire [31:0] _GEN_456; // @[FaultDetector.scala 177:34:@870.4]
  wire [3:0] _GEN_457; // @[FaultDetector.scala 177:34:@870.4]
  wire  _GEN_458; // @[FaultDetector.scala 177:34:@870.4]
  wire  reset_all_cpus; // @[FaultDetector.scala 485:28:@1142.4]
  wire  reset_all_cpus_out; // @[FaultDetector.scala 486:32:@1143.4]
  wire  reset_all_cpus_out_hold_clock; // @[FaultDetector.scala 487:39:@1144.4]
  wire  reset_all_cpus_out_hold_io_rst; // @[FaultDetector.scala 487:39:@1144.4]
  wire  reset_all_cpus_out_hold_io_o; // @[FaultDetector.scala 487:39:@1144.4]
  wire  reset_all_cpus_out_hold_io_i; // @[FaultDetector.scala 487:39:@1144.4]
  wire [1:0] _T_1946; // @[FaultDetector.scala 493:127:@1152.4]
  wire [2:0] _T_1947; // @[FaultDetector.scala 493:127:@1153.4]
  wire [2:0] _T_1948; // @[FaultDetector.scala 493:82:@1154.4]
  wire [2:0] _T_1949; // @[FaultDetector.scala 493:53:@1155.4]
  wire [2:0] _T_1950; // @[FaultDetector.scala 493:22:@1156.4]
  wire [2:0] _T_1959; // @[FaultDetector.scala 494:31:@1163.4]
  wire  _T_1969; // @[FaultDetector.scala 499:74:@1172.4]
  wire  _T_1971; // @[FaultDetector.scala 499:51:@1174.4]
  wire  _T_1972; // @[FaultDetector.scala 499:49:@1175.4]
  wire  _T_1974; // @[FaultDetector.scala 501:53:@1179.4]
  cpuRepair cpu_repair ( // @[FaultDetector.scala 394:26:@261.4]
    .clock(cpu_repair_clock),
    .reset(cpu_repair_reset),
    .io_fault(cpu_repair_io_fault),
    .io_cpus_ok(cpu_repair_io_cpus_ok),
    .io_reset_pending(cpu_repair_io_reset_pending),
    .io_ack_cpus_ok(cpu_repair_io_ack_cpus_ok),
    .io_stop_cpus(cpu_repair_io_stop_cpus),
    .io_latch_regs(cpu_repair_io_latch_regs),
    .io_reset_to_recovery(cpu_repair_io_reset_to_recovery),
    .io_reset_cpus(cpu_repair_io_reset_cpus),
    .io_reset_routing_logic(cpu_repair_io_reset_routing_logic),
    .io_cpu_in_interrupt(cpu_repair_io_cpu_in_interrupt)
  );
  signalHolder logic_reset_hold_0 ( // @[FaultDetector.scala 406:50:@276.4]
    .clock(logic_reset_hold_0_clock),
    .io_rst(logic_reset_hold_0_io_rst),
    .io_o(logic_reset_hold_0_io_o),
    .io_i(logic_reset_hold_0_io_i)
  );
  signalHolder logic_reset_hold_1 ( // @[FaultDetector.scala 406:87:@279.4]
    .clock(logic_reset_hold_1_clock),
    .io_rst(logic_reset_hold_1_io_rst),
    .io_o(logic_reset_hold_1_io_o),
    .io_i(logic_reset_hold_1_io_i)
  );
  signalHolder logic_reset_hold_2 ( // @[FaultDetector.scala 406:124:@282.4]
    .clock(logic_reset_hold_2_clock),
    .io_rst(logic_reset_hold_2_io_rst),
    .io_o(logic_reset_hold_2_io_o),
    .io_i(logic_reset_hold_2_io_i)
  );
  signalHolder cpu_reset_hold_0 ( // @[FaultDetector.scala 420:48:@303.4]
    .clock(cpu_reset_hold_0_clock),
    .io_rst(cpu_reset_hold_0_io_rst),
    .io_o(cpu_reset_hold_0_io_o),
    .io_i(cpu_reset_hold_0_io_i)
  );
  signalHolder cpu_reset_hold_1 ( // @[FaultDetector.scala 420:85:@306.4]
    .clock(cpu_reset_hold_1_clock),
    .io_rst(cpu_reset_hold_1_io_rst),
    .io_o(cpu_reset_hold_1_io_o),
    .io_i(cpu_reset_hold_1_io_i)
  );
  signalHolder cpu_reset_hold_2 ( // @[FaultDetector.scala 420:122:@309.4]
    .clock(cpu_reset_hold_2_clock),
    .io_rst(cpu_reset_hold_2_io_rst),
    .io_o(cpu_reset_hold_2_io_o),
    .io_i(cpu_reset_hold_2_io_i)
  );
  signalHolder reset_all_cpus_out_hold ( // @[FaultDetector.scala 487:39:@1144.4]
    .clock(reset_all_cpus_out_hold_clock),
    .io_rst(reset_all_cpus_out_hold_io_rst),
    .io_o(reset_all_cpus_out_hold_io_o),
    .io_i(reset_all_cpus_out_hold_io_i)
  );
  assign _T_397 = ~ reset_logic; // @[FaultDetector.scala 410:18:@286.4]
  assign _T_761 = {reset_routing_2,reset_routing_1}; // @[FaultDetector.scala 425:52:@321.4]
  assign _T_762 = {_T_761,reset_routing_0}; // @[FaultDetector.scala 425:52:@322.4]
  assign _T_764 = _T_762 != 3'h0; // @[FaultDetector.scala 425:59:@323.4]
  assign _T_1229 = io_cpu0_axi4_aw_valid != io_cpu1_axi4_aw_valid; // @[FaultDetector.scala 323:43:@326.4]
  assign _T_1230 = io_cpu0_axi4_w_valid != io_cpu1_axi4_w_valid; // @[FaultDetector.scala 324:42:@328.4]
  assign _T_1231 = io_cpu0_axi4_ar_valid != io_cpu1_axi4_ar_valid; // @[FaultDetector.scala 325:43:@330.4]
  assign _T_1232 = io_cpu0_axi4_b_ready != io_cpu1_axi4_b_ready; // @[FaultDetector.scala 327:42:@332.4]
  assign _T_1233 = io_cpu0_axi4_r_ready != io_cpu1_axi4_r_ready; // @[FaultDetector.scala 328:42:@334.4]
  assign _T_1234 = io_cpu0_axi4_aw_bits_id ^ io_cpu1_axi4_aw_bits_id; // @[FaultDetector.scala 330:46:@336.4]
  assign _T_1236 = _T_1234 != 4'h0; // @[FaultDetector.scala 330:67:@337.4]
  assign _T_1237 = io_cpu0_axi4_aw_bits_addr ^ io_cpu1_axi4_aw_bits_addr; // @[FaultDetector.scala 331:48:@339.4]
  assign _T_1239 = _T_1237 != 32'h0; // @[FaultDetector.scala 331:71:@340.4]
  assign _T_1240 = io_cpu0_axi4_aw_bits_len ^ io_cpu1_axi4_aw_bits_len; // @[FaultDetector.scala 332:47:@342.4]
  assign _T_1242 = _T_1240 != 8'h0; // @[FaultDetector.scala 332:69:@343.4]
  assign _T_1243 = io_cpu0_axi4_aw_bits_size ^ io_cpu1_axi4_aw_bits_size; // @[FaultDetector.scala 333:48:@345.4]
  assign _T_1245 = _T_1243 != 3'h0; // @[FaultDetector.scala 333:71:@346.4]
  assign _T_1246 = io_cpu0_axi4_aw_bits_burst ^ io_cpu1_axi4_aw_bits_burst; // @[FaultDetector.scala 334:49:@348.4]
  assign _T_1248 = _T_1246 != 2'h0; // @[FaultDetector.scala 334:73:@349.4]
  assign _T_1249 = io_cpu0_axi4_aw_bits_lock ^ io_cpu1_axi4_aw_bits_lock; // @[FaultDetector.scala 335:49:@351.4]
  assign _T_1252 = io_cpu0_axi4_aw_bits_cache ^ io_cpu1_axi4_aw_bits_cache; // @[FaultDetector.scala 336:50:@354.4]
  assign _T_1254 = _T_1252 != 4'h0; // @[FaultDetector.scala 336:74:@355.4]
  assign _T_1255 = io_cpu0_axi4_aw_bits_prot ^ io_cpu1_axi4_aw_bits_prot; // @[FaultDetector.scala 337:49:@357.4]
  assign _T_1257 = _T_1255 != 3'h0; // @[FaultDetector.scala 337:72:@358.4]
  assign _T_1258 = io_cpu0_axi4_aw_bits_qos ^ io_cpu1_axi4_aw_bits_qos; // @[FaultDetector.scala 338:48:@360.4]
  assign _T_1260 = _T_1258 != 4'h0; // @[FaultDetector.scala 338:70:@361.4]
  assign _T_1261 = io_cpu0_axi4_ar_bits_id ^ io_cpu1_axi4_ar_bits_id; // @[FaultDetector.scala 340:47:@363.4]
  assign _T_1263 = _T_1261 != 4'h0; // @[FaultDetector.scala 340:68:@364.4]
  assign _T_1264 = io_cpu0_axi4_ar_bits_addr ^ io_cpu1_axi4_ar_bits_addr; // @[FaultDetector.scala 341:49:@366.4]
  assign _T_1266 = _T_1264 != 32'h0; // @[FaultDetector.scala 341:72:@367.4]
  assign _T_1267 = io_cpu0_axi4_ar_bits_len ^ io_cpu1_axi4_ar_bits_len; // @[FaultDetector.scala 342:48:@369.4]
  assign _T_1269 = _T_1267 != 8'h0; // @[FaultDetector.scala 342:70:@370.4]
  assign _T_1270 = io_cpu0_axi4_ar_bits_size ^ io_cpu1_axi4_ar_bits_size; // @[FaultDetector.scala 343:49:@372.4]
  assign _T_1272 = _T_1270 != 3'h0; // @[FaultDetector.scala 343:72:@373.4]
  assign _T_1273 = io_cpu0_axi4_ar_bits_burst ^ io_cpu1_axi4_ar_bits_burst; // @[FaultDetector.scala 344:50:@375.4]
  assign _T_1275 = _T_1273 != 2'h0; // @[FaultDetector.scala 344:74:@376.4]
  assign _T_1276 = io_cpu0_axi4_ar_bits_lock ^ io_cpu1_axi4_ar_bits_lock; // @[FaultDetector.scala 345:49:@378.4]
  assign _T_1279 = io_cpu0_axi4_ar_bits_cache ^ io_cpu1_axi4_ar_bits_cache; // @[FaultDetector.scala 346:50:@381.4]
  assign _T_1281 = _T_1279 != 4'h0; // @[FaultDetector.scala 346:74:@382.4]
  assign _T_1282 = io_cpu0_axi4_ar_bits_prot ^ io_cpu1_axi4_ar_bits_prot; // @[FaultDetector.scala 347:49:@384.4]
  assign _T_1284 = _T_1282 != 3'h0; // @[FaultDetector.scala 347:72:@385.4]
  assign _T_1285 = io_cpu0_axi4_ar_bits_qos ^ io_cpu1_axi4_ar_bits_qos; // @[FaultDetector.scala 348:48:@387.4]
  assign _T_1287 = _T_1285 != 4'h0; // @[FaultDetector.scala 348:70:@388.4]
  assign _T_1288 = io_cpu0_axi4_w_bits_data ^ io_cpu1_axi4_w_bits_data; // @[FaultDetector.scala 350:48:@390.4]
  assign _T_1290 = _T_1288 != 32'h0; // @[FaultDetector.scala 350:70:@391.4]
  assign _T_1291 = io_cpu0_axi4_w_bits_strb ^ io_cpu1_axi4_w_bits_strb; // @[FaultDetector.scala 351:48:@393.4]
  assign _T_1293 = _T_1291 != 4'h0; // @[FaultDetector.scala 351:70:@394.4]
  assign _T_1294 = io_cpu0_axi4_w_bits_last ^ io_cpu1_axi4_w_bits_last; // @[FaultDetector.scala 352:48:@396.4]
  assign _T_1351 = _T_891_0_0 | _T_891_0_1; // @[FaultDetector.scala 354:46:@426.4]
  assign _T_1352 = _T_1351 | _T_891_0_2; // @[FaultDetector.scala 354:46:@427.4]
  assign _T_1353 = _T_1352 | _T_891_0_3; // @[FaultDetector.scala 354:46:@428.4]
  assign _T_1354 = _T_1353 | _T_891_0_4; // @[FaultDetector.scala 354:46:@429.4]
  assign _T_1355 = _T_1354 | _T_891_0_5; // @[FaultDetector.scala 354:46:@430.4]
  assign _T_1356 = _T_1355 | _T_891_0_6; // @[FaultDetector.scala 354:46:@431.4]
  assign _T_1357 = _T_1356 | _T_891_0_7; // @[FaultDetector.scala 354:46:@432.4]
  assign _T_1358 = _T_1357 | _T_891_0_8; // @[FaultDetector.scala 354:46:@433.4]
  assign _T_1359 = _T_1358 | _T_891_0_9; // @[FaultDetector.scala 354:46:@434.4]
  assign _T_1360 = _T_1359 | _T_891_0_10; // @[FaultDetector.scala 354:46:@435.4]
  assign _T_1361 = _T_1360 | _T_891_0_11; // @[FaultDetector.scala 354:46:@436.4]
  assign _T_1362 = _T_1361 | _T_891_0_12; // @[FaultDetector.scala 354:46:@437.4]
  assign _T_1363 = _T_1362 | _T_891_0_13; // @[FaultDetector.scala 354:46:@438.4]
  assign _T_1364 = _T_1363 | _T_891_0_14; // @[FaultDetector.scala 354:46:@439.4]
  assign _T_1365 = _T_1364 | _T_891_0_15; // @[FaultDetector.scala 354:46:@440.4]
  assign _T_1366 = _T_1365 | _T_891_0_16; // @[FaultDetector.scala 354:46:@441.4]
  assign _T_1367 = _T_1366 | _T_891_0_17; // @[FaultDetector.scala 354:46:@442.4]
  assign _T_1368 = _T_1367 | _T_891_0_18; // @[FaultDetector.scala 354:46:@443.4]
  assign _T_1369 = _T_1368 | _T_891_0_19; // @[FaultDetector.scala 354:46:@444.4]
  assign _T_1370 = _T_1369 | _T_891_0_20; // @[FaultDetector.scala 354:46:@445.4]
  assign _T_1371 = _T_1370 | _T_891_0_21; // @[FaultDetector.scala 354:46:@446.4]
  assign _T_1372 = _T_1371 | _T_891_0_22; // @[FaultDetector.scala 354:46:@447.4]
  assign _T_1373 = _T_1372 | _T_891_0_23; // @[FaultDetector.scala 354:46:@448.4]
  assign _T_1374 = _T_1373 | _T_891_0_24; // @[FaultDetector.scala 354:46:@449.4]
  assign _T_1375 = _T_1374 | _T_891_0_25; // @[FaultDetector.scala 354:46:@450.4]
  assign _T_1376 = io_cpu0_axi4_aw_valid != io_cpu2_axi4_aw_valid; // @[FaultDetector.scala 323:43:@452.4]
  assign _T_1377 = io_cpu0_axi4_w_valid != io_cpu2_axi4_w_valid; // @[FaultDetector.scala 324:42:@454.4]
  assign _T_1378 = io_cpu0_axi4_ar_valid != io_cpu2_axi4_ar_valid; // @[FaultDetector.scala 325:43:@456.4]
  assign _T_1379 = io_cpu0_axi4_b_ready != io_cpu2_axi4_b_ready; // @[FaultDetector.scala 327:42:@458.4]
  assign _T_1380 = io_cpu0_axi4_r_ready != io_cpu2_axi4_r_ready; // @[FaultDetector.scala 328:42:@460.4]
  assign _T_1381 = io_cpu0_axi4_aw_bits_id ^ io_cpu2_axi4_aw_bits_id; // @[FaultDetector.scala 330:46:@462.4]
  assign _T_1383 = _T_1381 != 4'h0; // @[FaultDetector.scala 330:67:@463.4]
  assign _T_1384 = io_cpu0_axi4_aw_bits_addr ^ io_cpu2_axi4_aw_bits_addr; // @[FaultDetector.scala 331:48:@465.4]
  assign _T_1386 = _T_1384 != 32'h0; // @[FaultDetector.scala 331:71:@466.4]
  assign _T_1387 = io_cpu0_axi4_aw_bits_len ^ io_cpu2_axi4_aw_bits_len; // @[FaultDetector.scala 332:47:@468.4]
  assign _T_1389 = _T_1387 != 8'h0; // @[FaultDetector.scala 332:69:@469.4]
  assign _T_1390 = io_cpu0_axi4_aw_bits_size ^ io_cpu2_axi4_aw_bits_size; // @[FaultDetector.scala 333:48:@471.4]
  assign _T_1392 = _T_1390 != 3'h0; // @[FaultDetector.scala 333:71:@472.4]
  assign _T_1393 = io_cpu0_axi4_aw_bits_burst ^ io_cpu2_axi4_aw_bits_burst; // @[FaultDetector.scala 334:49:@474.4]
  assign _T_1395 = _T_1393 != 2'h0; // @[FaultDetector.scala 334:73:@475.4]
  assign _T_1396 = io_cpu0_axi4_aw_bits_lock ^ io_cpu2_axi4_aw_bits_lock; // @[FaultDetector.scala 335:49:@477.4]
  assign _T_1399 = io_cpu0_axi4_aw_bits_cache ^ io_cpu2_axi4_aw_bits_cache; // @[FaultDetector.scala 336:50:@480.4]
  assign _T_1401 = _T_1399 != 4'h0; // @[FaultDetector.scala 336:74:@481.4]
  assign _T_1402 = io_cpu0_axi4_aw_bits_prot ^ io_cpu2_axi4_aw_bits_prot; // @[FaultDetector.scala 337:49:@483.4]
  assign _T_1404 = _T_1402 != 3'h0; // @[FaultDetector.scala 337:72:@484.4]
  assign _T_1405 = io_cpu0_axi4_aw_bits_qos ^ io_cpu2_axi4_aw_bits_qos; // @[FaultDetector.scala 338:48:@486.4]
  assign _T_1407 = _T_1405 != 4'h0; // @[FaultDetector.scala 338:70:@487.4]
  assign _T_1408 = io_cpu0_axi4_ar_bits_id ^ io_cpu2_axi4_ar_bits_id; // @[FaultDetector.scala 340:47:@489.4]
  assign _T_1410 = _T_1408 != 4'h0; // @[FaultDetector.scala 340:68:@490.4]
  assign _T_1411 = io_cpu0_axi4_ar_bits_addr ^ io_cpu2_axi4_ar_bits_addr; // @[FaultDetector.scala 341:49:@492.4]
  assign _T_1413 = _T_1411 != 32'h0; // @[FaultDetector.scala 341:72:@493.4]
  assign _T_1414 = io_cpu0_axi4_ar_bits_len ^ io_cpu2_axi4_ar_bits_len; // @[FaultDetector.scala 342:48:@495.4]
  assign _T_1416 = _T_1414 != 8'h0; // @[FaultDetector.scala 342:70:@496.4]
  assign _T_1417 = io_cpu0_axi4_ar_bits_size ^ io_cpu2_axi4_ar_bits_size; // @[FaultDetector.scala 343:49:@498.4]
  assign _T_1419 = _T_1417 != 3'h0; // @[FaultDetector.scala 343:72:@499.4]
  assign _T_1420 = io_cpu0_axi4_ar_bits_burst ^ io_cpu2_axi4_ar_bits_burst; // @[FaultDetector.scala 344:50:@501.4]
  assign _T_1422 = _T_1420 != 2'h0; // @[FaultDetector.scala 344:74:@502.4]
  assign _T_1423 = io_cpu0_axi4_ar_bits_lock ^ io_cpu2_axi4_ar_bits_lock; // @[FaultDetector.scala 345:49:@504.4]
  assign _T_1426 = io_cpu0_axi4_ar_bits_cache ^ io_cpu2_axi4_ar_bits_cache; // @[FaultDetector.scala 346:50:@507.4]
  assign _T_1428 = _T_1426 != 4'h0; // @[FaultDetector.scala 346:74:@508.4]
  assign _T_1429 = io_cpu0_axi4_ar_bits_prot ^ io_cpu2_axi4_ar_bits_prot; // @[FaultDetector.scala 347:49:@510.4]
  assign _T_1431 = _T_1429 != 3'h0; // @[FaultDetector.scala 347:72:@511.4]
  assign _T_1432 = io_cpu0_axi4_ar_bits_qos ^ io_cpu2_axi4_ar_bits_qos; // @[FaultDetector.scala 348:48:@513.4]
  assign _T_1434 = _T_1432 != 4'h0; // @[FaultDetector.scala 348:70:@514.4]
  assign _T_1435 = io_cpu0_axi4_w_bits_data ^ io_cpu2_axi4_w_bits_data; // @[FaultDetector.scala 350:48:@516.4]
  assign _T_1437 = _T_1435 != 32'h0; // @[FaultDetector.scala 350:70:@517.4]
  assign _T_1438 = io_cpu0_axi4_w_bits_strb ^ io_cpu2_axi4_w_bits_strb; // @[FaultDetector.scala 351:48:@519.4]
  assign _T_1440 = _T_1438 != 4'h0; // @[FaultDetector.scala 351:70:@520.4]
  assign _T_1441 = io_cpu0_axi4_w_bits_last ^ io_cpu2_axi4_w_bits_last; // @[FaultDetector.scala 352:48:@522.4]
  assign _T_1498 = _T_891_1_0 | _T_891_1_1; // @[FaultDetector.scala 354:46:@552.4]
  assign _T_1499 = _T_1498 | _T_891_1_2; // @[FaultDetector.scala 354:46:@553.4]
  assign _T_1500 = _T_1499 | _T_891_1_3; // @[FaultDetector.scala 354:46:@554.4]
  assign _T_1501 = _T_1500 | _T_891_1_4; // @[FaultDetector.scala 354:46:@555.4]
  assign _T_1502 = _T_1501 | _T_891_1_5; // @[FaultDetector.scala 354:46:@556.4]
  assign _T_1503 = _T_1502 | _T_891_1_6; // @[FaultDetector.scala 354:46:@557.4]
  assign _T_1504 = _T_1503 | _T_891_1_7; // @[FaultDetector.scala 354:46:@558.4]
  assign _T_1505 = _T_1504 | _T_891_1_8; // @[FaultDetector.scala 354:46:@559.4]
  assign _T_1506 = _T_1505 | _T_891_1_9; // @[FaultDetector.scala 354:46:@560.4]
  assign _T_1507 = _T_1506 | _T_891_1_10; // @[FaultDetector.scala 354:46:@561.4]
  assign _T_1508 = _T_1507 | _T_891_1_11; // @[FaultDetector.scala 354:46:@562.4]
  assign _T_1509 = _T_1508 | _T_891_1_12; // @[FaultDetector.scala 354:46:@563.4]
  assign _T_1510 = _T_1509 | _T_891_1_13; // @[FaultDetector.scala 354:46:@564.4]
  assign _T_1511 = _T_1510 | _T_891_1_14; // @[FaultDetector.scala 354:46:@565.4]
  assign _T_1512 = _T_1511 | _T_891_1_15; // @[FaultDetector.scala 354:46:@566.4]
  assign _T_1513 = _T_1512 | _T_891_1_16; // @[FaultDetector.scala 354:46:@567.4]
  assign _T_1514 = _T_1513 | _T_891_1_17; // @[FaultDetector.scala 354:46:@568.4]
  assign _T_1515 = _T_1514 | _T_891_1_18; // @[FaultDetector.scala 354:46:@569.4]
  assign _T_1516 = _T_1515 | _T_891_1_19; // @[FaultDetector.scala 354:46:@570.4]
  assign _T_1517 = _T_1516 | _T_891_1_20; // @[FaultDetector.scala 354:46:@571.4]
  assign _T_1518 = _T_1517 | _T_891_1_21; // @[FaultDetector.scala 354:46:@572.4]
  assign _T_1519 = _T_1518 | _T_891_1_22; // @[FaultDetector.scala 354:46:@573.4]
  assign _T_1520 = _T_1519 | _T_891_1_23; // @[FaultDetector.scala 354:46:@574.4]
  assign _T_1521 = _T_1520 | _T_891_1_24; // @[FaultDetector.scala 354:46:@575.4]
  assign _T_1522 = _T_1521 | _T_891_1_25; // @[FaultDetector.scala 354:46:@576.4]
  assign _T_1523 = io_cpu1_axi4_aw_valid != io_cpu2_axi4_aw_valid; // @[FaultDetector.scala 323:43:@578.4]
  assign _T_1524 = io_cpu1_axi4_w_valid != io_cpu2_axi4_w_valid; // @[FaultDetector.scala 324:42:@580.4]
  assign _T_1525 = io_cpu1_axi4_ar_valid != io_cpu2_axi4_ar_valid; // @[FaultDetector.scala 325:43:@582.4]
  assign _T_1526 = io_cpu1_axi4_b_ready != io_cpu2_axi4_b_ready; // @[FaultDetector.scala 327:42:@584.4]
  assign _T_1527 = io_cpu1_axi4_r_ready != io_cpu2_axi4_r_ready; // @[FaultDetector.scala 328:42:@586.4]
  assign _T_1528 = io_cpu1_axi4_aw_bits_id ^ io_cpu2_axi4_aw_bits_id; // @[FaultDetector.scala 330:46:@588.4]
  assign _T_1530 = _T_1528 != 4'h0; // @[FaultDetector.scala 330:67:@589.4]
  assign _T_1531 = io_cpu1_axi4_aw_bits_addr ^ io_cpu2_axi4_aw_bits_addr; // @[FaultDetector.scala 331:48:@591.4]
  assign _T_1533 = _T_1531 != 32'h0; // @[FaultDetector.scala 331:71:@592.4]
  assign _T_1534 = io_cpu1_axi4_aw_bits_len ^ io_cpu2_axi4_aw_bits_len; // @[FaultDetector.scala 332:47:@594.4]
  assign _T_1536 = _T_1534 != 8'h0; // @[FaultDetector.scala 332:69:@595.4]
  assign _T_1537 = io_cpu1_axi4_aw_bits_size ^ io_cpu2_axi4_aw_bits_size; // @[FaultDetector.scala 333:48:@597.4]
  assign _T_1539 = _T_1537 != 3'h0; // @[FaultDetector.scala 333:71:@598.4]
  assign _T_1540 = io_cpu1_axi4_aw_bits_burst ^ io_cpu2_axi4_aw_bits_burst; // @[FaultDetector.scala 334:49:@600.4]
  assign _T_1542 = _T_1540 != 2'h0; // @[FaultDetector.scala 334:73:@601.4]
  assign _T_1543 = io_cpu1_axi4_aw_bits_lock ^ io_cpu2_axi4_aw_bits_lock; // @[FaultDetector.scala 335:49:@603.4]
  assign _T_1546 = io_cpu1_axi4_aw_bits_cache ^ io_cpu2_axi4_aw_bits_cache; // @[FaultDetector.scala 336:50:@606.4]
  assign _T_1548 = _T_1546 != 4'h0; // @[FaultDetector.scala 336:74:@607.4]
  assign _T_1549 = io_cpu1_axi4_aw_bits_prot ^ io_cpu2_axi4_aw_bits_prot; // @[FaultDetector.scala 337:49:@609.4]
  assign _T_1551 = _T_1549 != 3'h0; // @[FaultDetector.scala 337:72:@610.4]
  assign _T_1552 = io_cpu1_axi4_aw_bits_qos ^ io_cpu2_axi4_aw_bits_qos; // @[FaultDetector.scala 338:48:@612.4]
  assign _T_1554 = _T_1552 != 4'h0; // @[FaultDetector.scala 338:70:@613.4]
  assign _T_1555 = io_cpu1_axi4_ar_bits_id ^ io_cpu2_axi4_ar_bits_id; // @[FaultDetector.scala 340:47:@615.4]
  assign _T_1557 = _T_1555 != 4'h0; // @[FaultDetector.scala 340:68:@616.4]
  assign _T_1558 = io_cpu1_axi4_ar_bits_addr ^ io_cpu2_axi4_ar_bits_addr; // @[FaultDetector.scala 341:49:@618.4]
  assign _T_1560 = _T_1558 != 32'h0; // @[FaultDetector.scala 341:72:@619.4]
  assign _T_1561 = io_cpu1_axi4_ar_bits_len ^ io_cpu2_axi4_ar_bits_len; // @[FaultDetector.scala 342:48:@621.4]
  assign _T_1563 = _T_1561 != 8'h0; // @[FaultDetector.scala 342:70:@622.4]
  assign _T_1564 = io_cpu1_axi4_ar_bits_size ^ io_cpu2_axi4_ar_bits_size; // @[FaultDetector.scala 343:49:@624.4]
  assign _T_1566 = _T_1564 != 3'h0; // @[FaultDetector.scala 343:72:@625.4]
  assign _T_1567 = io_cpu1_axi4_ar_bits_burst ^ io_cpu2_axi4_ar_bits_burst; // @[FaultDetector.scala 344:50:@627.4]
  assign _T_1569 = _T_1567 != 2'h0; // @[FaultDetector.scala 344:74:@628.4]
  assign _T_1570 = io_cpu1_axi4_ar_bits_lock ^ io_cpu2_axi4_ar_bits_lock; // @[FaultDetector.scala 345:49:@630.4]
  assign _T_1573 = io_cpu1_axi4_ar_bits_cache ^ io_cpu2_axi4_ar_bits_cache; // @[FaultDetector.scala 346:50:@633.4]
  assign _T_1575 = _T_1573 != 4'h0; // @[FaultDetector.scala 346:74:@634.4]
  assign _T_1576 = io_cpu1_axi4_ar_bits_prot ^ io_cpu2_axi4_ar_bits_prot; // @[FaultDetector.scala 347:49:@636.4]
  assign _T_1578 = _T_1576 != 3'h0; // @[FaultDetector.scala 347:72:@637.4]
  assign _T_1579 = io_cpu1_axi4_ar_bits_qos ^ io_cpu2_axi4_ar_bits_qos; // @[FaultDetector.scala 348:48:@639.4]
  assign _T_1581 = _T_1579 != 4'h0; // @[FaultDetector.scala 348:70:@640.4]
  assign _T_1582 = io_cpu1_axi4_w_bits_data ^ io_cpu2_axi4_w_bits_data; // @[FaultDetector.scala 350:48:@642.4]
  assign _T_1584 = _T_1582 != 32'h0; // @[FaultDetector.scala 350:70:@643.4]
  assign _T_1585 = io_cpu1_axi4_w_bits_strb ^ io_cpu2_axi4_w_bits_strb; // @[FaultDetector.scala 351:48:@645.4]
  assign _T_1587 = _T_1585 != 4'h0; // @[FaultDetector.scala 351:70:@646.4]
  assign _T_1588 = io_cpu1_axi4_w_bits_last ^ io_cpu2_axi4_w_bits_last; // @[FaultDetector.scala 352:48:@648.4]
  assign _T_1645 = _T_891_2_0 | _T_891_2_1; // @[FaultDetector.scala 354:46:@678.4]
  assign _T_1646 = _T_1645 | _T_891_2_2; // @[FaultDetector.scala 354:46:@679.4]
  assign _T_1647 = _T_1646 | _T_891_2_3; // @[FaultDetector.scala 354:46:@680.4]
  assign _T_1648 = _T_1647 | _T_891_2_4; // @[FaultDetector.scala 354:46:@681.4]
  assign _T_1649 = _T_1648 | _T_891_2_5; // @[FaultDetector.scala 354:46:@682.4]
  assign _T_1650 = _T_1649 | _T_891_2_6; // @[FaultDetector.scala 354:46:@683.4]
  assign _T_1651 = _T_1650 | _T_891_2_7; // @[FaultDetector.scala 354:46:@684.4]
  assign _T_1652 = _T_1651 | _T_891_2_8; // @[FaultDetector.scala 354:46:@685.4]
  assign _T_1653 = _T_1652 | _T_891_2_9; // @[FaultDetector.scala 354:46:@686.4]
  assign _T_1654 = _T_1653 | _T_891_2_10; // @[FaultDetector.scala 354:46:@687.4]
  assign _T_1655 = _T_1654 | _T_891_2_11; // @[FaultDetector.scala 354:46:@688.4]
  assign _T_1656 = _T_1655 | _T_891_2_12; // @[FaultDetector.scala 354:46:@689.4]
  assign _T_1657 = _T_1656 | _T_891_2_13; // @[FaultDetector.scala 354:46:@690.4]
  assign _T_1658 = _T_1657 | _T_891_2_14; // @[FaultDetector.scala 354:46:@691.4]
  assign _T_1659 = _T_1658 | _T_891_2_15; // @[FaultDetector.scala 354:46:@692.4]
  assign _T_1660 = _T_1659 | _T_891_2_16; // @[FaultDetector.scala 354:46:@693.4]
  assign _T_1661 = _T_1660 | _T_891_2_17; // @[FaultDetector.scala 354:46:@694.4]
  assign _T_1662 = _T_1661 | _T_891_2_18; // @[FaultDetector.scala 354:46:@695.4]
  assign _T_1663 = _T_1662 | _T_891_2_19; // @[FaultDetector.scala 354:46:@696.4]
  assign _T_1664 = _T_1663 | _T_891_2_20; // @[FaultDetector.scala 354:46:@697.4]
  assign _T_1665 = _T_1664 | _T_891_2_21; // @[FaultDetector.scala 354:46:@698.4]
  assign _T_1666 = _T_1665 | _T_891_2_22; // @[FaultDetector.scala 354:46:@699.4]
  assign _T_1667 = _T_1666 | _T_891_2_23; // @[FaultDetector.scala 354:46:@700.4]
  assign _T_1668 = _T_1667 | _T_891_2_24; // @[FaultDetector.scala 354:46:@701.4]
  assign _T_1669 = _T_1668 | _T_891_2_25; // @[FaultDetector.scala 354:46:@702.4]
  assign _T_1672 = {1'h0,_T_768_0}; // @[Cat.scala 30:58:@704.4]
  assign _T_1673 = {_T_1672,_T_768_1}; // @[Cat.scala 30:58:@705.4]
  assign _T_1674 = {_T_1673,_T_768_2}; // @[Cat.scala 30:58:@706.4]
  assign invalid = _T_764 ? 4'h0 : _T_1674; // @[FaultDetector.scala 358:8:@707.4]
  assign _GEN_0 = reset_logic ? 1'h1 : reset_logic_reg; // @[FaultDetector.scala 434:28:@714.4]
  assign _GEN_5 = reset_logic ? 3'h0 : invalid_reg; // @[FaultDetector.scala 434:28:@714.4]
  assign _T_1693 = invalid == 4'h0; // @[FaultDetector.scala 444:18:@724.6]
  assign _GEN_7 = _T_1693 ? 1'h0 : _GEN_0; // @[FaultDetector.scala 444:27:@725.6]
  assign _GEN_8 = _T_1693 ? 1'h1 : cpu_back_online_reg; // @[FaultDetector.scala 444:27:@725.6]
  assign _GEN_9 = reset_logic_reg ? _GEN_7 : _GEN_0; // @[FaultDetector.scala 443:25:@723.4]
  assign _GEN_10 = reset_logic_reg ? _GEN_8 : cpu_back_online_reg; // @[FaultDetector.scala 443:25:@723.4]
  assign _GEN_11 = ack_back_online ? 1'h0 : _GEN_10; // @[FaultDetector.scala 450:25:@730.4]
  assign _T_1698 = invalid != 4'h0; // @[FaultDetector.scala 456:16:@734.4]
  assign _T_1701 = reset_logic_reg == 1'h0; // @[FaultDetector.scala 456:27:@736.4]
  assign _T_1702 = _T_1698 & _T_1701; // @[FaultDetector.scala 456:24:@737.4]
  assign _GEN_12 = _T_1702 ? invalid : {{1'd0}, _GEN_5}; // @[FaultDetector.scala 456:52:@738.4]
  assign _T_1704 = invalid_reg != 3'h0; // @[FaultDetector.scala 460:20:@741.4]
  assign _T_1705 = ~ invalid_reg; // @[FaultDetector.scala 462:21:@743.6]
  assign _GEN_13 = _T_1704 ? _T_1705 : 3'h0; // @[FaultDetector.scala 460:29:@742.4]
  assign _T_1709 = cpu_reset_im[0]; // @[FaultDetector.scala 473:30:@753.4]
  assign _T_1710 = cpu_reset_im[1]; // @[FaultDetector.scala 473:30:@757.4]
  assign _T_1711 = cpu_reset_im[2]; // @[FaultDetector.scala 473:30:@761.4]
  assign invalid_bool_0 = faulty_cpu[0]; // @[FaultDetector.scala 477:33:@764.4]
  assign invalid_bool_1 = faulty_cpu[1]; // @[FaultDetector.scala 477:33:@765.4]
  assign invalid_bool_2 = faulty_cpu[2]; // @[FaultDetector.scala 477:33:@766.4]
  assign _T_1713 = reset_routing_0 == 1'h0; // @[FaultDetector.scala 121:8:@767.4]
  assign _GEN_15 = invalid_bool_0 ? 1'h0 : _T_429_aw_ready; // @[FaultDetector.scala 125:21:@772.6]
  assign _GEN_16 = invalid_bool_0 ? 1'h0 : _T_429_w_ready; // @[FaultDetector.scala 125:21:@772.6]
  assign _GEN_17 = invalid_bool_0 ? 1'h0 : _T_429_ar_ready; // @[FaultDetector.scala 125:21:@772.6]
  assign _GEN_18 = invalid_bool_0 ? 1'h0 : _T_429_b_valid; // @[FaultDetector.scala 125:21:@772.6]
  assign _GEN_19 = invalid_bool_0 ? 4'h0 : _T_429_b_bits_id; // @[FaultDetector.scala 125:21:@772.6]
  assign _GEN_20 = invalid_bool_0 ? 2'h0 : _T_429_b_bits_resp; // @[FaultDetector.scala 125:21:@772.6]
  assign _GEN_21 = invalid_bool_0 ? 1'h0 : _T_429_r_valid; // @[FaultDetector.scala 125:21:@772.6]
  assign _GEN_22 = invalid_bool_0 ? 4'h0 : _T_429_r_bits_id; // @[FaultDetector.scala 125:21:@772.6]
  assign _GEN_23 = invalid_bool_0 ? 2'h0 : _T_429_r_bits_resp; // @[FaultDetector.scala 125:21:@772.6]
  assign _GEN_24 = invalid_bool_0 ? 1'h0 : _T_429_r_bits_last; // @[FaultDetector.scala 125:21:@772.6]
  assign _GEN_25 = invalid_bool_0 ? 32'h0 : _T_429_r_bits_data; // @[FaultDetector.scala 125:21:@772.6]
  assign _GEN_26 = _T_1713 ? _GEN_15 : _T_429_aw_ready; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_37 = _T_1713 ? _GEN_16 : _T_429_w_ready; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_43 = _T_1713 ? _GEN_18 : _T_429_b_valid; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_44 = _T_1713 ? _GEN_19 : _T_429_b_bits_id; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_45 = _T_1713 ? _GEN_20 : _T_429_b_bits_resp; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_46 = _T_1713 ? _GEN_17 : _T_429_ar_ready; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_58 = _T_1713 ? _GEN_21 : _T_429_r_valid; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_59 = _T_1713 ? _GEN_22 : _T_429_r_bits_id; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_60 = _T_1713 ? _GEN_25 : _T_429_r_bits_data; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_61 = _T_1713 ? _GEN_23 : _T_429_r_bits_resp; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_62 = _T_1713 ? _GEN_24 : _T_429_r_bits_last; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_63 = _T_1713 ? _T_487_aw_ready : _T_429_aw_ready; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_64 = _T_1713 ? _T_429_aw_valid : _T_487_aw_valid; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_65 = _T_1713 ? _T_429_aw_bits_id : _T_487_aw_bits_id; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_66 = _T_1713 ? _T_429_aw_bits_addr : _T_487_aw_bits_addr; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_67 = _T_1713 ? _T_429_aw_bits_len : _T_487_aw_bits_len; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_68 = _T_1713 ? _T_429_aw_bits_size : _T_487_aw_bits_size; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_69 = _T_1713 ? _T_429_aw_bits_burst : _T_487_aw_bits_burst; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_70 = _T_1713 ? _T_429_aw_bits_lock : _T_487_aw_bits_lock; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_71 = _T_1713 ? _T_429_aw_bits_cache : _T_487_aw_bits_cache; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_72 = _T_1713 ? _T_429_aw_bits_prot : _T_487_aw_bits_prot; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_73 = _T_1713 ? _T_429_aw_bits_qos : _T_487_aw_bits_qos; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_74 = _T_1713 ? _T_487_w_ready : _T_429_w_ready; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_75 = _T_1713 ? _T_429_w_valid : _T_487_w_valid; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_76 = _T_1713 ? _T_429_w_bits_data : _T_487_w_bits_data; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_77 = _T_1713 ? _T_429_w_bits_strb : _T_487_w_bits_strb; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_78 = _T_1713 ? _T_429_w_bits_last : _T_487_w_bits_last; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_79 = _T_1713 ? _T_429_b_ready : _T_487_b_ready; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_80 = _T_1713 ? _T_487_b_valid : _T_429_b_valid; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_81 = _T_1713 ? _T_487_b_bits_id : _T_429_b_bits_id; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_82 = _T_1713 ? _T_487_b_bits_resp : _T_429_b_bits_resp; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_83 = _T_1713 ? _T_487_ar_ready : _T_429_ar_ready; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_84 = _T_1713 ? _T_429_ar_valid : _T_487_ar_valid; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_85 = _T_1713 ? _T_429_ar_bits_id : _T_487_ar_bits_id; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_86 = _T_1713 ? _T_429_ar_bits_addr : _T_487_ar_bits_addr; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_87 = _T_1713 ? _T_429_ar_bits_len : _T_487_ar_bits_len; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_88 = _T_1713 ? _T_429_ar_bits_size : _T_487_ar_bits_size; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_89 = _T_1713 ? _T_429_ar_bits_burst : _T_487_ar_bits_burst; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_90 = _T_1713 ? _T_429_ar_bits_lock : _T_487_ar_bits_lock; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_91 = _T_1713 ? _T_429_ar_bits_cache : _T_487_ar_bits_cache; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_92 = _T_1713 ? _T_429_ar_bits_prot : _T_487_ar_bits_prot; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_93 = _T_1713 ? _T_429_ar_bits_qos : _T_487_ar_bits_qos; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_94 = _T_1713 ? _T_429_r_ready : _T_487_r_ready; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_95 = _T_1713 ? _T_487_r_valid : _T_429_r_valid; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_96 = _T_1713 ? _T_487_r_bits_id : _T_429_r_bits_id; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_97 = _T_1713 ? _T_487_r_bits_data : _T_429_r_bits_data; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_98 = _T_1713 ? _T_487_r_bits_resp : _T_429_r_bits_resp; // @[FaultDetector.scala 121:15:@768.4]
  assign _GEN_99 = _T_1713 ? _T_487_r_bits_last : _T_429_r_bits_last; // @[FaultDetector.scala 121:15:@768.4]
  assign _T_1726 = reset_routing_1 == 1'h0; // @[FaultDetector.scala 121:8:@790.4]
  assign _GEN_137 = invalid_bool_1 ? 1'h0 : _T_545_aw_ready; // @[FaultDetector.scala 125:21:@795.6]
  assign _GEN_138 = invalid_bool_1 ? 1'h0 : _T_545_w_ready; // @[FaultDetector.scala 125:21:@795.6]
  assign _GEN_139 = invalid_bool_1 ? 1'h0 : _T_545_ar_ready; // @[FaultDetector.scala 125:21:@795.6]
  assign _GEN_140 = invalid_bool_1 ? 1'h0 : _T_545_b_valid; // @[FaultDetector.scala 125:21:@795.6]
  assign _GEN_141 = invalid_bool_1 ? 4'h0 : _T_545_b_bits_id; // @[FaultDetector.scala 125:21:@795.6]
  assign _GEN_142 = invalid_bool_1 ? 2'h0 : _T_545_b_bits_resp; // @[FaultDetector.scala 125:21:@795.6]
  assign _GEN_143 = invalid_bool_1 ? 1'h0 : _T_545_r_valid; // @[FaultDetector.scala 125:21:@795.6]
  assign _GEN_144 = invalid_bool_1 ? 4'h0 : _T_545_r_bits_id; // @[FaultDetector.scala 125:21:@795.6]
  assign _GEN_145 = invalid_bool_1 ? 2'h0 : _T_545_r_bits_resp; // @[FaultDetector.scala 125:21:@795.6]
  assign _GEN_146 = invalid_bool_1 ? 1'h0 : _T_545_r_bits_last; // @[FaultDetector.scala 125:21:@795.6]
  assign _GEN_147 = invalid_bool_1 ? 32'h0 : _T_545_r_bits_data; // @[FaultDetector.scala 125:21:@795.6]
  assign _GEN_148 = _T_1726 ? _GEN_137 : _T_545_aw_ready; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_159 = _T_1726 ? _GEN_138 : _T_545_w_ready; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_165 = _T_1726 ? _GEN_140 : _T_545_b_valid; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_166 = _T_1726 ? _GEN_141 : _T_545_b_bits_id; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_167 = _T_1726 ? _GEN_142 : _T_545_b_bits_resp; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_168 = _T_1726 ? _GEN_139 : _T_545_ar_ready; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_180 = _T_1726 ? _GEN_143 : _T_545_r_valid; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_181 = _T_1726 ? _GEN_144 : _T_545_r_bits_id; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_182 = _T_1726 ? _GEN_147 : _T_545_r_bits_data; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_183 = _T_1726 ? _GEN_145 : _T_545_r_bits_resp; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_184 = _T_1726 ? _GEN_146 : _T_545_r_bits_last; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_185 = _T_1726 ? _T_603_aw_ready : _T_545_aw_ready; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_186 = _T_1726 ? _T_545_aw_valid : _T_603_aw_valid; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_187 = _T_1726 ? _T_545_aw_bits_id : _T_603_aw_bits_id; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_188 = _T_1726 ? _T_545_aw_bits_addr : _T_603_aw_bits_addr; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_189 = _T_1726 ? _T_545_aw_bits_len : _T_603_aw_bits_len; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_190 = _T_1726 ? _T_545_aw_bits_size : _T_603_aw_bits_size; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_191 = _T_1726 ? _T_545_aw_bits_burst : _T_603_aw_bits_burst; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_192 = _T_1726 ? _T_545_aw_bits_lock : _T_603_aw_bits_lock; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_193 = _T_1726 ? _T_545_aw_bits_cache : _T_603_aw_bits_cache; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_194 = _T_1726 ? _T_545_aw_bits_prot : _T_603_aw_bits_prot; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_195 = _T_1726 ? _T_545_aw_bits_qos : _T_603_aw_bits_qos; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_196 = _T_1726 ? _T_603_w_ready : _T_545_w_ready; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_197 = _T_1726 ? _T_545_w_valid : _T_603_w_valid; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_198 = _T_1726 ? _T_545_w_bits_data : _T_603_w_bits_data; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_199 = _T_1726 ? _T_545_w_bits_strb : _T_603_w_bits_strb; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_200 = _T_1726 ? _T_545_w_bits_last : _T_603_w_bits_last; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_201 = _T_1726 ? _T_545_b_ready : _T_603_b_ready; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_202 = _T_1726 ? _T_603_b_valid : _T_545_b_valid; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_203 = _T_1726 ? _T_603_b_bits_id : _T_545_b_bits_id; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_204 = _T_1726 ? _T_603_b_bits_resp : _T_545_b_bits_resp; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_205 = _T_1726 ? _T_603_ar_ready : _T_545_ar_ready; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_206 = _T_1726 ? _T_545_ar_valid : _T_603_ar_valid; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_207 = _T_1726 ? _T_545_ar_bits_id : _T_603_ar_bits_id; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_208 = _T_1726 ? _T_545_ar_bits_addr : _T_603_ar_bits_addr; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_209 = _T_1726 ? _T_545_ar_bits_len : _T_603_ar_bits_len; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_210 = _T_1726 ? _T_545_ar_bits_size : _T_603_ar_bits_size; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_211 = _T_1726 ? _T_545_ar_bits_burst : _T_603_ar_bits_burst; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_212 = _T_1726 ? _T_545_ar_bits_lock : _T_603_ar_bits_lock; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_213 = _T_1726 ? _T_545_ar_bits_cache : _T_603_ar_bits_cache; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_214 = _T_1726 ? _T_545_ar_bits_prot : _T_603_ar_bits_prot; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_215 = _T_1726 ? _T_545_ar_bits_qos : _T_603_ar_bits_qos; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_216 = _T_1726 ? _T_545_r_ready : _T_603_r_ready; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_217 = _T_1726 ? _T_603_r_valid : _T_545_r_valid; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_218 = _T_1726 ? _T_603_r_bits_id : _T_545_r_bits_id; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_219 = _T_1726 ? _T_603_r_bits_data : _T_545_r_bits_data; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_220 = _T_1726 ? _T_603_r_bits_resp : _T_545_r_bits_resp; // @[FaultDetector.scala 121:15:@791.4]
  assign _GEN_221 = _T_1726 ? _T_603_r_bits_last : _T_545_r_bits_last; // @[FaultDetector.scala 121:15:@791.4]
  assign _T_1739 = reset_routing_2 == 1'h0; // @[FaultDetector.scala 121:8:@813.4]
  assign _GEN_259 = invalid_bool_2 ? 1'h0 : _T_661_aw_ready; // @[FaultDetector.scala 125:21:@818.6]
  assign _GEN_260 = invalid_bool_2 ? 1'h0 : _T_661_w_ready; // @[FaultDetector.scala 125:21:@818.6]
  assign _GEN_261 = invalid_bool_2 ? 1'h0 : _T_661_ar_ready; // @[FaultDetector.scala 125:21:@818.6]
  assign _GEN_262 = invalid_bool_2 ? 1'h0 : _T_661_b_valid; // @[FaultDetector.scala 125:21:@818.6]
  assign _GEN_263 = invalid_bool_2 ? 4'h0 : _T_661_b_bits_id; // @[FaultDetector.scala 125:21:@818.6]
  assign _GEN_264 = invalid_bool_2 ? 2'h0 : _T_661_b_bits_resp; // @[FaultDetector.scala 125:21:@818.6]
  assign _GEN_265 = invalid_bool_2 ? 1'h0 : _T_661_r_valid; // @[FaultDetector.scala 125:21:@818.6]
  assign _GEN_266 = invalid_bool_2 ? 4'h0 : _T_661_r_bits_id; // @[FaultDetector.scala 125:21:@818.6]
  assign _GEN_267 = invalid_bool_2 ? 2'h0 : _T_661_r_bits_resp; // @[FaultDetector.scala 125:21:@818.6]
  assign _GEN_268 = invalid_bool_2 ? 1'h0 : _T_661_r_bits_last; // @[FaultDetector.scala 125:21:@818.6]
  assign _GEN_269 = invalid_bool_2 ? 32'h0 : _T_661_r_bits_data; // @[FaultDetector.scala 125:21:@818.6]
  assign _GEN_270 = _T_1739 ? _GEN_259 : _T_661_aw_ready; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_281 = _T_1739 ? _GEN_260 : _T_661_w_ready; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_287 = _T_1739 ? _GEN_262 : _T_661_b_valid; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_288 = _T_1739 ? _GEN_263 : _T_661_b_bits_id; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_289 = _T_1739 ? _GEN_264 : _T_661_b_bits_resp; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_290 = _T_1739 ? _GEN_261 : _T_661_ar_ready; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_302 = _T_1739 ? _GEN_265 : _T_661_r_valid; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_303 = _T_1739 ? _GEN_266 : _T_661_r_bits_id; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_304 = _T_1739 ? _GEN_269 : _T_661_r_bits_data; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_305 = _T_1739 ? _GEN_267 : _T_661_r_bits_resp; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_306 = _T_1739 ? _GEN_268 : _T_661_r_bits_last; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_307 = _T_1739 ? _T_719_aw_ready : _T_661_aw_ready; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_308 = _T_1739 ? _T_661_aw_valid : _T_719_aw_valid; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_309 = _T_1739 ? _T_661_aw_bits_id : _T_719_aw_bits_id; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_310 = _T_1739 ? _T_661_aw_bits_addr : _T_719_aw_bits_addr; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_311 = _T_1739 ? _T_661_aw_bits_len : _T_719_aw_bits_len; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_312 = _T_1739 ? _T_661_aw_bits_size : _T_719_aw_bits_size; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_313 = _T_1739 ? _T_661_aw_bits_burst : _T_719_aw_bits_burst; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_314 = _T_1739 ? _T_661_aw_bits_lock : _T_719_aw_bits_lock; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_315 = _T_1739 ? _T_661_aw_bits_cache : _T_719_aw_bits_cache; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_316 = _T_1739 ? _T_661_aw_bits_prot : _T_719_aw_bits_prot; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_317 = _T_1739 ? _T_661_aw_bits_qos : _T_719_aw_bits_qos; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_318 = _T_1739 ? _T_719_w_ready : _T_661_w_ready; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_319 = _T_1739 ? _T_661_w_valid : _T_719_w_valid; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_320 = _T_1739 ? _T_661_w_bits_data : _T_719_w_bits_data; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_321 = _T_1739 ? _T_661_w_bits_strb : _T_719_w_bits_strb; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_322 = _T_1739 ? _T_661_w_bits_last : _T_719_w_bits_last; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_323 = _T_1739 ? _T_661_b_ready : _T_719_b_ready; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_324 = _T_1739 ? _T_719_b_valid : _T_661_b_valid; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_325 = _T_1739 ? _T_719_b_bits_id : _T_661_b_bits_id; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_326 = _T_1739 ? _T_719_b_bits_resp : _T_661_b_bits_resp; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_327 = _T_1739 ? _T_719_ar_ready : _T_661_ar_ready; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_328 = _T_1739 ? _T_661_ar_valid : _T_719_ar_valid; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_329 = _T_1739 ? _T_661_ar_bits_id : _T_719_ar_bits_id; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_330 = _T_1739 ? _T_661_ar_bits_addr : _T_719_ar_bits_addr; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_331 = _T_1739 ? _T_661_ar_bits_len : _T_719_ar_bits_len; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_332 = _T_1739 ? _T_661_ar_bits_size : _T_719_ar_bits_size; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_333 = _T_1739 ? _T_661_ar_bits_burst : _T_719_ar_bits_burst; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_334 = _T_1739 ? _T_661_ar_bits_lock : _T_719_ar_bits_lock; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_335 = _T_1739 ? _T_661_ar_bits_cache : _T_719_ar_bits_cache; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_336 = _T_1739 ? _T_661_ar_bits_prot : _T_719_ar_bits_prot; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_337 = _T_1739 ? _T_661_ar_bits_qos : _T_719_ar_bits_qos; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_338 = _T_1739 ? _T_661_r_ready : _T_719_r_ready; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_339 = _T_1739 ? _T_719_r_valid : _T_661_r_valid; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_340 = _T_1739 ? _T_719_r_bits_id : _T_661_r_bits_id; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_341 = _T_1739 ? _T_719_r_bits_data : _T_661_r_bits_data; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_342 = _T_1739 ? _T_719_r_bits_resp : _T_661_r_bits_resp; // @[FaultDetector.scala 121:15:@814.4]
  assign _GEN_343 = _T_1739 ? _T_719_r_bits_last : _T_661_r_bits_last; // @[FaultDetector.scala 121:15:@814.4]
  assign _T_1752 = invalid_reg == 3'h6; // @[FaultDetector.scala 177:24:@869.4]
  assign _T_1753 = axiBusInternal1_aw_valid | axiBusInternal2_aw_valid; // @[FaultDetector.scala 179:56:@871.6]
  assign _T_1754 = axiBusInternal1_w_valid | axiBusInternal2_w_valid; // @[FaultDetector.scala 180:56:@873.6]
  assign _T_1755 = axiBusInternal1_ar_valid | axiBusInternal2_ar_valid; // @[FaultDetector.scala 181:56:@875.6]
  assign _T_1756 = axiBusInternal1_b_ready | axiBusInternal2_b_ready; // @[FaultDetector.scala 183:54:@877.6]
  assign _T_1757 = axiBusInternal1_r_ready | axiBusInternal2_r_ready; // @[FaultDetector.scala 184:54:@879.6]
  assign _T_1758 = axiBusInternal1_aw_bits_id | axiBusInternal2_aw_bits_id; // @[FaultDetector.scala 186:66:@881.6]
  assign _T_1759 = axiBusInternal1_aw_bits_addr | axiBusInternal2_aw_bits_addr; // @[FaultDetector.scala 187:66:@883.6]
  assign _T_1760 = axiBusInternal1_aw_bits_len | axiBusInternal2_aw_bits_len; // @[FaultDetector.scala 188:66:@885.6]
  assign _T_1761 = axiBusInternal1_aw_bits_size | axiBusInternal2_aw_bits_size; // @[FaultDetector.scala 189:66:@887.6]
  assign _T_1762 = axiBusInternal1_aw_bits_burst | axiBusInternal2_aw_bits_burst; // @[FaultDetector.scala 190:66:@889.6]
  assign _T_1763 = axiBusInternal1_aw_bits_lock | axiBusInternal2_aw_bits_lock; // @[FaultDetector.scala 191:66:@891.6]
  assign _T_1764 = axiBusInternal1_aw_bits_cache | axiBusInternal2_aw_bits_cache; // @[FaultDetector.scala 192:66:@893.6]
  assign _T_1765 = axiBusInternal1_aw_bits_prot | axiBusInternal2_aw_bits_prot; // @[FaultDetector.scala 193:66:@895.6]
  assign _T_1766 = axiBusInternal1_aw_bits_qos | axiBusInternal2_aw_bits_qos; // @[FaultDetector.scala 194:66:@897.6]
  assign _T_1767 = axiBusInternal1_ar_bits_id | axiBusInternal2_ar_bits_id; // @[FaultDetector.scala 196:66:@899.6]
  assign _T_1768 = axiBusInternal1_ar_bits_addr | axiBusInternal2_ar_bits_addr; // @[FaultDetector.scala 197:66:@901.6]
  assign _T_1769 = axiBusInternal1_ar_bits_len | axiBusInternal2_ar_bits_len; // @[FaultDetector.scala 198:66:@903.6]
  assign _T_1770 = axiBusInternal1_ar_bits_size | axiBusInternal2_ar_bits_size; // @[FaultDetector.scala 199:66:@905.6]
  assign _T_1771 = axiBusInternal1_ar_bits_burst | axiBusInternal2_ar_bits_burst; // @[FaultDetector.scala 200:66:@907.6]
  assign _T_1772 = axiBusInternal1_ar_bits_lock | axiBusInternal2_ar_bits_lock; // @[FaultDetector.scala 201:66:@909.6]
  assign _T_1773 = axiBusInternal1_ar_bits_cache | axiBusInternal2_ar_bits_cache; // @[FaultDetector.scala 202:66:@911.6]
  assign _T_1774 = axiBusInternal1_ar_bits_prot | axiBusInternal2_ar_bits_prot; // @[FaultDetector.scala 203:66:@913.6]
  assign _T_1775 = axiBusInternal1_ar_bits_qos | axiBusInternal2_ar_bits_qos; // @[FaultDetector.scala 204:66:@915.6]
  assign _T_1776 = axiBusInternal1_w_bits_data | axiBusInternal2_w_bits_data; // @[FaultDetector.scala 206:62:@917.6]
  assign _T_1777 = axiBusInternal1_w_bits_strb | axiBusInternal2_w_bits_strb; // @[FaultDetector.scala 207:62:@919.6]
  assign _T_1778 = axiBusInternal1_w_bits_last | axiBusInternal2_w_bits_last; // @[FaultDetector.scala 208:62:@921.6]
  assign _T_1780 = invalid_reg == 3'h5; // @[FaultDetector.scala 210:30:@925.6]
  assign _T_1781 = axiBusInternal0_aw_valid | axiBusInternal2_aw_valid; // @[FaultDetector.scala 212:56:@927.8]
  assign _T_1782 = axiBusInternal0_w_valid | axiBusInternal2_w_valid; // @[FaultDetector.scala 213:56:@929.8]
  assign _T_1783 = axiBusInternal0_ar_valid | axiBusInternal2_ar_valid; // @[FaultDetector.scala 214:56:@931.8]
  assign _T_1784 = axiBusInternal0_b_ready | axiBusInternal2_b_ready; // @[FaultDetector.scala 216:54:@933.8]
  assign _T_1785 = axiBusInternal0_r_ready | axiBusInternal2_r_ready; // @[FaultDetector.scala 217:54:@935.8]
  assign _T_1786 = axiBusInternal0_aw_bits_id | axiBusInternal2_aw_bits_id; // @[FaultDetector.scala 219:66:@937.8]
  assign _T_1787 = axiBusInternal0_aw_bits_addr | axiBusInternal2_aw_bits_addr; // @[FaultDetector.scala 220:66:@939.8]
  assign _T_1788 = axiBusInternal0_aw_bits_len | axiBusInternal2_aw_bits_len; // @[FaultDetector.scala 221:66:@941.8]
  assign _T_1789 = axiBusInternal0_aw_bits_size | axiBusInternal2_aw_bits_size; // @[FaultDetector.scala 222:66:@943.8]
  assign _T_1790 = axiBusInternal0_aw_bits_burst | axiBusInternal2_aw_bits_burst; // @[FaultDetector.scala 223:66:@945.8]
  assign _T_1791 = axiBusInternal0_aw_bits_lock | axiBusInternal2_aw_bits_lock; // @[FaultDetector.scala 224:66:@947.8]
  assign _T_1792 = axiBusInternal0_aw_bits_cache | axiBusInternal2_aw_bits_cache; // @[FaultDetector.scala 225:66:@949.8]
  assign _T_1793 = axiBusInternal0_aw_bits_prot | axiBusInternal2_aw_bits_prot; // @[FaultDetector.scala 226:66:@951.8]
  assign _T_1794 = axiBusInternal0_aw_bits_qos | axiBusInternal2_aw_bits_qos; // @[FaultDetector.scala 227:66:@953.8]
  assign _T_1795 = axiBusInternal0_ar_bits_id | axiBusInternal2_ar_bits_id; // @[FaultDetector.scala 229:66:@955.8]
  assign _T_1796 = axiBusInternal0_ar_bits_addr | axiBusInternal2_ar_bits_addr; // @[FaultDetector.scala 230:66:@957.8]
  assign _T_1797 = axiBusInternal0_ar_bits_len | axiBusInternal2_ar_bits_len; // @[FaultDetector.scala 231:66:@959.8]
  assign _T_1798 = axiBusInternal0_ar_bits_size | axiBusInternal2_ar_bits_size; // @[FaultDetector.scala 232:66:@961.8]
  assign _T_1799 = axiBusInternal0_ar_bits_burst | axiBusInternal2_ar_bits_burst; // @[FaultDetector.scala 233:66:@963.8]
  assign _T_1800 = axiBusInternal0_ar_bits_lock | axiBusInternal2_ar_bits_lock; // @[FaultDetector.scala 234:66:@965.8]
  assign _T_1801 = axiBusInternal0_ar_bits_cache | axiBusInternal2_ar_bits_cache; // @[FaultDetector.scala 235:66:@967.8]
  assign _T_1802 = axiBusInternal0_ar_bits_prot | axiBusInternal2_ar_bits_prot; // @[FaultDetector.scala 236:66:@969.8]
  assign _T_1803 = axiBusInternal0_ar_bits_qos | axiBusInternal2_ar_bits_qos; // @[FaultDetector.scala 237:66:@971.8]
  assign _T_1804 = axiBusInternal0_w_bits_data | axiBusInternal2_w_bits_data; // @[FaultDetector.scala 239:62:@973.8]
  assign _T_1805 = axiBusInternal0_w_bits_strb | axiBusInternal2_w_bits_strb; // @[FaultDetector.scala 240:62:@975.8]
  assign _T_1806 = axiBusInternal0_w_bits_last | axiBusInternal2_w_bits_last; // @[FaultDetector.scala 241:62:@977.8]
  assign _T_1808 = invalid_reg == 3'h3; // @[FaultDetector.scala 243:30:@981.8]
  assign _T_1809 = axiBusInternal0_aw_valid | axiBusInternal1_aw_valid; // @[FaultDetector.scala 245:56:@983.10]
  assign _T_1810 = axiBusInternal0_w_valid | axiBusInternal1_w_valid; // @[FaultDetector.scala 246:56:@985.10]
  assign _T_1811 = axiBusInternal0_ar_valid | axiBusInternal1_ar_valid; // @[FaultDetector.scala 247:56:@987.10]
  assign _T_1812 = axiBusInternal0_b_ready | axiBusInternal1_b_ready; // @[FaultDetector.scala 249:54:@989.10]
  assign _T_1813 = axiBusInternal0_r_ready | axiBusInternal1_r_ready; // @[FaultDetector.scala 250:54:@991.10]
  assign _T_1814 = axiBusInternal0_aw_bits_id | axiBusInternal1_aw_bits_id; // @[FaultDetector.scala 252:66:@993.10]
  assign _T_1815 = axiBusInternal0_aw_bits_addr | axiBusInternal1_aw_bits_addr; // @[FaultDetector.scala 253:66:@995.10]
  assign _T_1816 = axiBusInternal0_aw_bits_len | axiBusInternal1_aw_bits_len; // @[FaultDetector.scala 254:66:@997.10]
  assign _T_1817 = axiBusInternal0_aw_bits_size | axiBusInternal1_aw_bits_size; // @[FaultDetector.scala 255:66:@999.10]
  assign _T_1818 = axiBusInternal0_aw_bits_burst | axiBusInternal1_aw_bits_burst; // @[FaultDetector.scala 256:66:@1001.10]
  assign _T_1819 = axiBusInternal0_aw_bits_lock | axiBusInternal1_aw_bits_lock; // @[FaultDetector.scala 257:66:@1003.10]
  assign _T_1820 = axiBusInternal0_aw_bits_cache | axiBusInternal1_aw_bits_cache; // @[FaultDetector.scala 258:66:@1005.10]
  assign _T_1821 = axiBusInternal0_aw_bits_prot | axiBusInternal1_aw_bits_prot; // @[FaultDetector.scala 259:66:@1007.10]
  assign _T_1822 = axiBusInternal0_aw_bits_qos | axiBusInternal1_aw_bits_qos; // @[FaultDetector.scala 260:66:@1009.10]
  assign _T_1823 = axiBusInternal0_ar_bits_id | axiBusInternal1_ar_bits_id; // @[FaultDetector.scala 262:66:@1011.10]
  assign _T_1824 = axiBusInternal0_ar_bits_addr | axiBusInternal1_ar_bits_addr; // @[FaultDetector.scala 263:66:@1013.10]
  assign _T_1825 = axiBusInternal0_ar_bits_len | axiBusInternal1_ar_bits_len; // @[FaultDetector.scala 264:66:@1015.10]
  assign _T_1826 = axiBusInternal0_ar_bits_size | axiBusInternal1_ar_bits_size; // @[FaultDetector.scala 265:66:@1017.10]
  assign _T_1827 = axiBusInternal0_ar_bits_burst | axiBusInternal1_ar_bits_burst; // @[FaultDetector.scala 266:66:@1019.10]
  assign _T_1828 = axiBusInternal0_ar_bits_lock | axiBusInternal1_ar_bits_lock; // @[FaultDetector.scala 267:66:@1021.10]
  assign _T_1829 = axiBusInternal0_ar_bits_cache | axiBusInternal1_ar_bits_cache; // @[FaultDetector.scala 268:66:@1023.10]
  assign _T_1830 = axiBusInternal0_ar_bits_prot | axiBusInternal1_ar_bits_prot; // @[FaultDetector.scala 269:66:@1025.10]
  assign _T_1831 = axiBusInternal0_ar_bits_qos | axiBusInternal1_ar_bits_qos; // @[FaultDetector.scala 270:66:@1027.10]
  assign _T_1832 = axiBusInternal0_w_bits_data | axiBusInternal1_w_bits_data; // @[FaultDetector.scala 272:62:@1029.10]
  assign _T_1833 = axiBusInternal0_w_bits_strb | axiBusInternal1_w_bits_strb; // @[FaultDetector.scala 273:62:@1031.10]
  assign _T_1834 = axiBusInternal0_w_bits_last | axiBusInternal1_w_bits_last; // @[FaultDetector.scala 274:62:@1033.10]
  assign _T_1838 = _T_1809 | axiBusInternal2_aw_valid; // @[FaultDetector.scala 279:80:@1039.10]
  assign _T_1842 = _T_1810 | axiBusInternal2_w_valid; // @[FaultDetector.scala 280:80:@1043.10]
  assign _T_1846 = _T_1811 | axiBusInternal2_ar_valid; // @[FaultDetector.scala 281:80:@1047.10]
  assign _T_1850 = _T_1812 | axiBusInternal2_b_ready; // @[FaultDetector.scala 283:79:@1051.10]
  assign _T_1854 = _T_1813 | axiBusInternal2_r_ready; // @[FaultDetector.scala 284:79:@1055.10]
  assign _T_1858 = _T_1814 | axiBusInternal2_aw_bits_id; // @[FaultDetector.scala 286:81:@1059.10]
  assign _T_1862 = _T_1815 | axiBusInternal2_aw_bits_addr; // @[FaultDetector.scala 287:81:@1063.10]
  assign _T_1866 = _T_1816 | axiBusInternal2_aw_bits_len; // @[FaultDetector.scala 288:81:@1067.10]
  assign _T_1870 = _T_1817 | axiBusInternal2_aw_bits_size; // @[FaultDetector.scala 289:81:@1071.10]
  assign _T_1874 = _T_1818 | axiBusInternal2_aw_bits_burst; // @[FaultDetector.scala 290:81:@1075.10]
  assign _T_1878 = _T_1819 | axiBusInternal2_aw_bits_lock; // @[FaultDetector.scala 291:81:@1079.10]
  assign _T_1882 = _T_1820 | axiBusInternal2_aw_bits_cache; // @[FaultDetector.scala 292:81:@1083.10]
  assign _T_1886 = _T_1821 | axiBusInternal2_aw_bits_prot; // @[FaultDetector.scala 293:81:@1087.10]
  assign _T_1890 = _T_1822 | axiBusInternal2_aw_bits_qos; // @[FaultDetector.scala 294:81:@1091.10]
  assign _T_1894 = _T_1823 | axiBusInternal2_ar_bits_id; // @[FaultDetector.scala 296:81:@1095.10]
  assign _T_1898 = _T_1824 | axiBusInternal2_ar_bits_addr; // @[FaultDetector.scala 297:81:@1099.10]
  assign _T_1902 = _T_1825 | axiBusInternal2_ar_bits_len; // @[FaultDetector.scala 298:81:@1103.10]
  assign _T_1906 = _T_1826 | axiBusInternal2_ar_bits_size; // @[FaultDetector.scala 299:81:@1107.10]
  assign _T_1910 = _T_1827 | axiBusInternal2_ar_bits_burst; // @[FaultDetector.scala 300:81:@1111.10]
  assign _T_1914 = _T_1828 | axiBusInternal2_ar_bits_lock; // @[FaultDetector.scala 301:81:@1115.10]
  assign _T_1918 = _T_1829 | axiBusInternal2_ar_bits_cache; // @[FaultDetector.scala 302:81:@1119.10]
  assign _T_1922 = _T_1830 | axiBusInternal2_ar_bits_prot; // @[FaultDetector.scala 303:81:@1123.10]
  assign _T_1926 = _T_1831 | axiBusInternal2_ar_bits_qos; // @[FaultDetector.scala 304:81:@1127.10]
  assign _T_1930 = _T_1832 | axiBusInternal2_w_bits_data; // @[FaultDetector.scala 306:79:@1131.10]
  assign _T_1934 = _T_1833 | axiBusInternal2_w_bits_strb; // @[FaultDetector.scala 307:79:@1135.10]
  assign _T_1938 = _T_1834 | axiBusInternal2_w_bits_last; // @[FaultDetector.scala 308:79:@1139.10]
  assign _GEN_381 = _T_1808 ? _T_1809 : _T_1838; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_382 = _T_1808 ? _T_1810 : _T_1842; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_383 = _T_1808 ? _T_1811 : _T_1846; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_384 = _T_1808 ? _T_1812 : _T_1850; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_385 = _T_1808 ? _T_1813 : _T_1854; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_386 = _T_1808 ? _T_1814 : _T_1858; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_387 = _T_1808 ? _T_1815 : _T_1862; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_388 = _T_1808 ? _T_1816 : _T_1866; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_389 = _T_1808 ? _T_1817 : _T_1870; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_390 = _T_1808 ? _T_1818 : _T_1874; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_391 = _T_1808 ? _T_1819 : _T_1878; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_392 = _T_1808 ? _T_1820 : _T_1882; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_393 = _T_1808 ? _T_1821 : _T_1886; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_394 = _T_1808 ? _T_1822 : _T_1890; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_395 = _T_1808 ? _T_1823 : _T_1894; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_396 = _T_1808 ? _T_1824 : _T_1898; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_397 = _T_1808 ? _T_1825 : _T_1902; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_398 = _T_1808 ? _T_1826 : _T_1906; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_399 = _T_1808 ? _T_1827 : _T_1910; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_400 = _T_1808 ? _T_1828 : _T_1914; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_401 = _T_1808 ? _T_1829 : _T_1918; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_402 = _T_1808 ? _T_1830 : _T_1922; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_403 = _T_1808 ? _T_1831 : _T_1926; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_404 = _T_1808 ? _T_1832 : _T_1930; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_405 = _T_1808 ? _T_1833 : _T_1934; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_406 = _T_1808 ? _T_1834 : _T_1938; // @[FaultDetector.scala 243:40:@982.8]
  assign _GEN_407 = _T_1780 ? _T_1781 : _GEN_381; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_408 = _T_1780 ? _T_1782 : _GEN_382; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_409 = _T_1780 ? _T_1783 : _GEN_383; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_410 = _T_1780 ? _T_1784 : _GEN_384; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_411 = _T_1780 ? _T_1785 : _GEN_385; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_412 = _T_1780 ? _T_1786 : _GEN_386; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_413 = _T_1780 ? _T_1787 : _GEN_387; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_414 = _T_1780 ? _T_1788 : _GEN_388; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_415 = _T_1780 ? _T_1789 : _GEN_389; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_416 = _T_1780 ? _T_1790 : _GEN_390; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_417 = _T_1780 ? _T_1791 : _GEN_391; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_418 = _T_1780 ? _T_1792 : _GEN_392; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_419 = _T_1780 ? _T_1793 : _GEN_393; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_420 = _T_1780 ? _T_1794 : _GEN_394; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_421 = _T_1780 ? _T_1795 : _GEN_395; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_422 = _T_1780 ? _T_1796 : _GEN_396; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_423 = _T_1780 ? _T_1797 : _GEN_397; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_424 = _T_1780 ? _T_1798 : _GEN_398; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_425 = _T_1780 ? _T_1799 : _GEN_399; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_426 = _T_1780 ? _T_1800 : _GEN_400; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_427 = _T_1780 ? _T_1801 : _GEN_401; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_428 = _T_1780 ? _T_1802 : _GEN_402; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_429 = _T_1780 ? _T_1803 : _GEN_403; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_430 = _T_1780 ? _T_1804 : _GEN_404; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_431 = _T_1780 ? _T_1805 : _GEN_405; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_432 = _T_1780 ? _T_1806 : _GEN_406; // @[FaultDetector.scala 210:40:@926.6]
  assign _GEN_433 = _T_1752 ? _T_1753 : _GEN_407; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_434 = _T_1752 ? _T_1754 : _GEN_408; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_435 = _T_1752 ? _T_1755 : _GEN_409; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_436 = _T_1752 ? _T_1756 : _GEN_410; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_437 = _T_1752 ? _T_1757 : _GEN_411; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_438 = _T_1752 ? _T_1758 : _GEN_412; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_439 = _T_1752 ? _T_1759 : _GEN_413; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_440 = _T_1752 ? _T_1760 : _GEN_414; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_441 = _T_1752 ? _T_1761 : _GEN_415; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_442 = _T_1752 ? _T_1762 : _GEN_416; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_443 = _T_1752 ? _T_1763 : _GEN_417; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_444 = _T_1752 ? _T_1764 : _GEN_418; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_445 = _T_1752 ? _T_1765 : _GEN_419; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_446 = _T_1752 ? _T_1766 : _GEN_420; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_447 = _T_1752 ? _T_1767 : _GEN_421; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_448 = _T_1752 ? _T_1768 : _GEN_422; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_449 = _T_1752 ? _T_1769 : _GEN_423; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_450 = _T_1752 ? _T_1770 : _GEN_424; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_451 = _T_1752 ? _T_1771 : _GEN_425; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_452 = _T_1752 ? _T_1772 : _GEN_426; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_453 = _T_1752 ? _T_1773 : _GEN_427; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_454 = _T_1752 ? _T_1774 : _GEN_428; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_455 = _T_1752 ? _T_1775 : _GEN_429; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_456 = _T_1752 ? _T_1776 : _GEN_430; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_457 = _T_1752 ? _T_1777 : _GEN_431; // @[FaultDetector.scala 177:34:@870.4]
  assign _GEN_458 = _T_1752 ? _T_1778 : _GEN_432; // @[FaultDetector.scala 177:34:@870.4]
  assign _T_1946 = {cpu_reset_out_2,cpu_reset_out_1}; // @[FaultDetector.scala 493:127:@1152.4]
  assign _T_1947 = {_T_1946,cpu_reset_out_0}; // @[FaultDetector.scala 493:127:@1153.4]
  assign _T_1948 = io_disable_reset ? 3'h0 : _T_1947; // @[FaultDetector.scala 493:82:@1154.4]
  assign _T_1949 = reset_logic ? 3'h0 : _T_1948; // @[FaultDetector.scala 493:53:@1155.4]
  assign _T_1950 = reset_all_cpus_out ? 3'h7 : _T_1949; // @[FaultDetector.scala 493:22:@1156.4]
  assign _T_1959 = reset_logic ? 3'h0 : _GEN_13; // @[FaultDetector.scala 494:31:@1163.4]
  assign _T_1969 = _T_1947 != 3'h0; // @[FaultDetector.scala 499:74:@1172.4]
  assign _T_1971 = ~ _T_1969; // @[FaultDetector.scala 499:51:@1174.4]
  assign _T_1972 = _T_1704 & _T_1971; // @[FaultDetector.scala 499:49:@1175.4]
  assign _T_1974 = reset_all_cpus_out | io_cpu_reset_feedback; // @[FaultDetector.scala 501:53:@1179.4]
  assign io_invalid = _GEN_5;
  assign io_cpu0_axi4_aw_ready = _GEN_26;
  assign io_cpu0_axi4_w_ready = _GEN_37;
  assign io_cpu0_axi4_b_valid = _GEN_43;
  assign io_cpu0_axi4_b_bits_id = _GEN_44;
  assign io_cpu0_axi4_b_bits_resp = _GEN_45;
  assign io_cpu0_axi4_ar_ready = _GEN_46;
  assign io_cpu0_axi4_r_valid = _GEN_58;
  assign io_cpu0_axi4_r_bits_id = _GEN_59;
  assign io_cpu0_axi4_r_bits_data = _GEN_60;
  assign io_cpu0_axi4_r_bits_resp = _GEN_61;
  assign io_cpu0_axi4_r_bits_last = _GEN_62;
  assign io_cpu1_axi4_aw_ready = _GEN_148;
  assign io_cpu1_axi4_w_ready = _GEN_159;
  assign io_cpu1_axi4_b_valid = _GEN_165;
  assign io_cpu1_axi4_b_bits_id = _GEN_166;
  assign io_cpu1_axi4_b_bits_resp = _GEN_167;
  assign io_cpu1_axi4_ar_ready = _GEN_168;
  assign io_cpu1_axi4_r_valid = _GEN_180;
  assign io_cpu1_axi4_r_bits_id = _GEN_181;
  assign io_cpu1_axi4_r_bits_data = _GEN_182;
  assign io_cpu1_axi4_r_bits_resp = _GEN_183;
  assign io_cpu1_axi4_r_bits_last = _GEN_184;
  assign io_cpu2_axi4_aw_ready = _GEN_270;
  assign io_cpu2_axi4_w_ready = _GEN_281;
  assign io_cpu2_axi4_b_valid = _GEN_287;
  assign io_cpu2_axi4_b_bits_id = _GEN_288;
  assign io_cpu2_axi4_b_bits_resp = _GEN_289;
  assign io_cpu2_axi4_ar_ready = _GEN_290;
  assign io_cpu2_axi4_r_valid = _GEN_302;
  assign io_cpu2_axi4_r_bits_id = _GEN_303;
  assign io_cpu2_axi4_r_bits_data = _GEN_304;
  assign io_cpu2_axi4_r_bits_resp = _GEN_305;
  assign io_cpu2_axi4_r_bits_last = _GEN_306;
  assign io_out_axi4_aw_valid = _GEN_433;
  assign io_out_axi4_aw_bits_id = _GEN_438;
  assign io_out_axi4_aw_bits_addr = _GEN_439;
  assign io_out_axi4_aw_bits_len = _GEN_440;
  assign io_out_axi4_aw_bits_size = _GEN_441;
  assign io_out_axi4_aw_bits_burst = _GEN_442;
  assign io_out_axi4_aw_bits_lock = _GEN_443;
  assign io_out_axi4_aw_bits_cache = _GEN_444;
  assign io_out_axi4_aw_bits_prot = _GEN_445;
  assign io_out_axi4_aw_bits_qos = _GEN_446;
  assign io_out_axi4_w_valid = _GEN_434;
  assign io_out_axi4_w_bits_data = _GEN_456;
  assign io_out_axi4_w_bits_strb = _GEN_457;
  assign io_out_axi4_w_bits_last = _GEN_458;
  assign io_out_axi4_b_ready = _GEN_436;
  assign io_out_axi4_ar_valid = _GEN_435;
  assign io_out_axi4_ar_bits_id = _GEN_447;
  assign io_out_axi4_ar_bits_addr = _GEN_448;
  assign io_out_axi4_ar_bits_len = _GEN_449;
  assign io_out_axi4_ar_bits_size = _GEN_450;
  assign io_out_axi4_ar_bits_burst = _GEN_451;
  assign io_out_axi4_ar_bits_lock = _GEN_452;
  assign io_out_axi4_ar_bits_cache = _GEN_453;
  assign io_out_axi4_ar_bits_prot = _GEN_454;
  assign io_out_axi4_ar_bits_qos = _GEN_455;
  assign io_out_axi4_r_ready = _GEN_437;
  assign io_fault_reset_vector = _T_1959;
  assign io_reset_cpu = _T_1950;
  assign io_stop_all_cpus = cpu_repair_io_stop_cpus;
  assign io_latch_registers = cpu_repair_io_latch_regs;
  assign io_reset_to_recovery = cpu_repair_io_reset_to_recovery;
  assign io_cpu_back_online = cpu_back_online_reg;
  assign cpu_repair_clock = clock;
  assign cpu_repair_reset = reset;
  assign axiBusInternal0_aw_ready = io_out_axi4_aw_ready;
  assign axiBusInternal0_aw_valid = _T_487_aw_valid;
  assign axiBusInternal0_aw_bits_id = _T_487_aw_bits_id;
  assign axiBusInternal0_aw_bits_addr = _T_487_aw_bits_addr;
  assign axiBusInternal0_aw_bits_len = _T_487_aw_bits_len;
  assign axiBusInternal0_aw_bits_size = _T_487_aw_bits_size;
  assign axiBusInternal0_aw_bits_burst = _T_487_aw_bits_burst;
  assign axiBusInternal0_aw_bits_lock = _T_487_aw_bits_lock;
  assign axiBusInternal0_aw_bits_cache = _T_487_aw_bits_cache;
  assign axiBusInternal0_aw_bits_prot = _T_487_aw_bits_prot;
  assign axiBusInternal0_aw_bits_qos = _T_487_aw_bits_qos;
  assign axiBusInternal0_w_ready = io_out_axi4_w_ready;
  assign axiBusInternal0_w_valid = _T_487_w_valid;
  assign axiBusInternal0_w_bits_data = _T_487_w_bits_data;
  assign axiBusInternal0_w_bits_strb = _T_487_w_bits_strb;
  assign axiBusInternal0_w_bits_last = _T_487_w_bits_last;
  assign axiBusInternal0_b_ready = _T_487_b_ready;
  assign axiBusInternal0_b_valid = io_out_axi4_b_valid;
  assign axiBusInternal0_b_bits_id = io_out_axi4_b_bits_id;
  assign axiBusInternal0_b_bits_resp = io_out_axi4_b_bits_resp;
  assign axiBusInternal0_ar_ready = io_out_axi4_ar_ready;
  assign axiBusInternal0_ar_valid = _T_487_ar_valid;
  assign axiBusInternal0_ar_bits_id = _T_487_ar_bits_id;
  assign axiBusInternal0_ar_bits_addr = _T_487_ar_bits_addr;
  assign axiBusInternal0_ar_bits_len = _T_487_ar_bits_len;
  assign axiBusInternal0_ar_bits_size = _T_487_ar_bits_size;
  assign axiBusInternal0_ar_bits_burst = _T_487_ar_bits_burst;
  assign axiBusInternal0_ar_bits_lock = _T_487_ar_bits_lock;
  assign axiBusInternal0_ar_bits_cache = _T_487_ar_bits_cache;
  assign axiBusInternal0_ar_bits_prot = _T_487_ar_bits_prot;
  assign axiBusInternal0_ar_bits_qos = _T_487_ar_bits_qos;
  assign axiBusInternal0_r_ready = _T_487_r_ready;
  assign axiBusInternal0_r_valid = io_out_axi4_r_valid;
  assign axiBusInternal0_r_bits_id = io_out_axi4_r_bits_id;
  assign axiBusInternal0_r_bits_data = io_out_axi4_r_bits_data;
  assign axiBusInternal0_r_bits_resp = io_out_axi4_r_bits_resp;
  assign axiBusInternal0_r_bits_last = io_out_axi4_r_bits_last;
  assign axiBusInternal1_aw_ready = io_out_axi4_aw_ready;
  assign axiBusInternal1_aw_valid = _T_603_aw_valid;
  assign axiBusInternal1_aw_bits_id = _T_603_aw_bits_id;
  assign axiBusInternal1_aw_bits_addr = _T_603_aw_bits_addr;
  assign axiBusInternal1_aw_bits_len = _T_603_aw_bits_len;
  assign axiBusInternal1_aw_bits_size = _T_603_aw_bits_size;
  assign axiBusInternal1_aw_bits_burst = _T_603_aw_bits_burst;
  assign axiBusInternal1_aw_bits_lock = _T_603_aw_bits_lock;
  assign axiBusInternal1_aw_bits_cache = _T_603_aw_bits_cache;
  assign axiBusInternal1_aw_bits_prot = _T_603_aw_bits_prot;
  assign axiBusInternal1_aw_bits_qos = _T_603_aw_bits_qos;
  assign axiBusInternal1_w_ready = io_out_axi4_w_ready;
  assign axiBusInternal1_w_valid = _T_603_w_valid;
  assign axiBusInternal1_w_bits_data = _T_603_w_bits_data;
  assign axiBusInternal1_w_bits_strb = _T_603_w_bits_strb;
  assign axiBusInternal1_w_bits_last = _T_603_w_bits_last;
  assign axiBusInternal1_b_ready = _T_603_b_ready;
  assign axiBusInternal1_b_valid = io_out_axi4_b_valid;
  assign axiBusInternal1_b_bits_id = io_out_axi4_b_bits_id;
  assign axiBusInternal1_b_bits_resp = io_out_axi4_b_bits_resp;
  assign axiBusInternal1_ar_ready = io_out_axi4_ar_ready;
  assign axiBusInternal1_ar_valid = _T_603_ar_valid;
  assign axiBusInternal1_ar_bits_id = _T_603_ar_bits_id;
  assign axiBusInternal1_ar_bits_addr = _T_603_ar_bits_addr;
  assign axiBusInternal1_ar_bits_len = _T_603_ar_bits_len;
  assign axiBusInternal1_ar_bits_size = _T_603_ar_bits_size;
  assign axiBusInternal1_ar_bits_burst = _T_603_ar_bits_burst;
  assign axiBusInternal1_ar_bits_lock = _T_603_ar_bits_lock;
  assign axiBusInternal1_ar_bits_cache = _T_603_ar_bits_cache;
  assign axiBusInternal1_ar_bits_prot = _T_603_ar_bits_prot;
  assign axiBusInternal1_ar_bits_qos = _T_603_ar_bits_qos;
  assign axiBusInternal1_r_ready = _T_603_r_ready;
  assign axiBusInternal1_r_valid = io_out_axi4_r_valid;
  assign axiBusInternal1_r_bits_id = io_out_axi4_r_bits_id;
  assign axiBusInternal1_r_bits_data = io_out_axi4_r_bits_data;
  assign axiBusInternal1_r_bits_resp = io_out_axi4_r_bits_resp;
  assign axiBusInternal1_r_bits_last = io_out_axi4_r_bits_last;
  assign axiBusInternal2_aw_ready = io_out_axi4_aw_ready;
  assign axiBusInternal2_aw_valid = _T_719_aw_valid;
  assign axiBusInternal2_aw_bits_id = _T_719_aw_bits_id;
  assign axiBusInternal2_aw_bits_addr = _T_719_aw_bits_addr;
  assign axiBusInternal2_aw_bits_len = _T_719_aw_bits_len;
  assign axiBusInternal2_aw_bits_size = _T_719_aw_bits_size;
  assign axiBusInternal2_aw_bits_burst = _T_719_aw_bits_burst;
  assign axiBusInternal2_aw_bits_lock = _T_719_aw_bits_lock;
  assign axiBusInternal2_aw_bits_cache = _T_719_aw_bits_cache;
  assign axiBusInternal2_aw_bits_prot = _T_719_aw_bits_prot;
  assign axiBusInternal2_aw_bits_qos = _T_719_aw_bits_qos;
  assign axiBusInternal2_w_ready = io_out_axi4_w_ready;
  assign axiBusInternal2_w_valid = _T_719_w_valid;
  assign axiBusInternal2_w_bits_data = _T_719_w_bits_data;
  assign axiBusInternal2_w_bits_strb = _T_719_w_bits_strb;
  assign axiBusInternal2_w_bits_last = _T_719_w_bits_last;
  assign axiBusInternal2_b_ready = _T_719_b_ready;
  assign axiBusInternal2_b_valid = io_out_axi4_b_valid;
  assign axiBusInternal2_b_bits_id = io_out_axi4_b_bits_id;
  assign axiBusInternal2_b_bits_resp = io_out_axi4_b_bits_resp;
  assign axiBusInternal2_ar_ready = io_out_axi4_ar_ready;
  assign axiBusInternal2_ar_valid = _T_719_ar_valid;
  assign axiBusInternal2_ar_bits_id = _T_719_ar_bits_id;
  assign axiBusInternal2_ar_bits_addr = _T_719_ar_bits_addr;
  assign axiBusInternal2_ar_bits_len = _T_719_ar_bits_len;
  assign axiBusInternal2_ar_bits_size = _T_719_ar_bits_size;
  assign axiBusInternal2_ar_bits_burst = _T_719_ar_bits_burst;
  assign axiBusInternal2_ar_bits_lock = _T_719_ar_bits_lock;
  assign axiBusInternal2_ar_bits_cache = _T_719_ar_bits_cache;
  assign axiBusInternal2_ar_bits_prot = _T_719_ar_bits_prot;
  assign axiBusInternal2_ar_bits_qos = _T_719_ar_bits_qos;
  assign axiBusInternal2_r_ready = _T_719_r_ready;
  assign axiBusInternal2_r_valid = io_out_axi4_r_valid;
  assign axiBusInternal2_r_bits_id = io_out_axi4_r_bits_id;
  assign axiBusInternal2_r_bits_data = io_out_axi4_r_bits_data;
  assign axiBusInternal2_r_bits_resp = io_out_axi4_r_bits_resp;
  assign axiBusInternal2_r_bits_last = io_out_axi4_r_bits_last;
  assign reset_logic = cpu_repair_io_reset_routing_logic;
  assign reset_routing_0 = logic_reset_hold_0_io_o;
  assign reset_routing_1 = logic_reset_hold_1_io_o;
  assign reset_routing_2 = logic_reset_hold_2_io_o;
  assign logic_reset_hold_0_clock = clock;
  assign logic_reset_hold_1_clock = clock;
  assign logic_reset_hold_2_clock = clock;
  assign logic_reset_hold_0_io_rst = reset_logic;
  assign logic_reset_hold_0_io_i = _T_397;
  assign logic_reset_hold_1_io_rst = reset_logic;
  assign logic_reset_hold_1_io_i = _T_397;
  assign logic_reset_hold_2_io_rst = reset_logic;
  assign logic_reset_hold_2_io_i = _T_397;
  assign cpu_reset_hold_0_clock = clock;
  assign cpu_reset_hold_1_clock = clock;
  assign cpu_reset_hold_2_clock = clock;
  assign cpu_reset_out_0 = cpu_reset_hold_0_io_o;
  assign cpu_reset_out_1 = cpu_reset_hold_1_io_o;
  assign cpu_reset_out_2 = cpu_reset_hold_2_io_o;
  assign _T_768_0 = _T_1375;
  assign _T_768_1 = _T_1522;
  assign _T_768_2 = _T_1669;
  assign _T_891_0_0 = _T_1229;
  assign _T_891_0_1 = _T_1230;
  assign _T_891_0_2 = _T_1231;
  assign _T_891_0_3 = _T_1232;
  assign _T_891_0_4 = _T_1233;
  assign _T_891_0_5 = _T_1236;
  assign _T_891_0_6 = _T_1239;
  assign _T_891_0_7 = _T_1242;
  assign _T_891_0_8 = _T_1245;
  assign _T_891_0_9 = _T_1248;
  assign _T_891_0_10 = _T_1249;
  assign _T_891_0_11 = _T_1254;
  assign _T_891_0_12 = _T_1257;
  assign _T_891_0_13 = _T_1260;
  assign _T_891_0_14 = _T_1263;
  assign _T_891_0_15 = _T_1266;
  assign _T_891_0_16 = _T_1269;
  assign _T_891_0_17 = _T_1272;
  assign _T_891_0_18 = _T_1275;
  assign _T_891_0_19 = _T_1276;
  assign _T_891_0_20 = _T_1281;
  assign _T_891_0_21 = _T_1284;
  assign _T_891_0_22 = _T_1287;
  assign _T_891_0_23 = _T_1290;
  assign _T_891_0_24 = _T_1293;
  assign _T_891_0_25 = _T_1294;
  assign _T_891_1_0 = _T_1376;
  assign _T_891_1_1 = _T_1377;
  assign _T_891_1_2 = _T_1378;
  assign _T_891_1_3 = _T_1379;
  assign _T_891_1_4 = _T_1380;
  assign _T_891_1_5 = _T_1383;
  assign _T_891_1_6 = _T_1386;
  assign _T_891_1_7 = _T_1389;
  assign _T_891_1_8 = _T_1392;
  assign _T_891_1_9 = _T_1395;
  assign _T_891_1_10 = _T_1396;
  assign _T_891_1_11 = _T_1401;
  assign _T_891_1_12 = _T_1404;
  assign _T_891_1_13 = _T_1407;
  assign _T_891_1_14 = _T_1410;
  assign _T_891_1_15 = _T_1413;
  assign _T_891_1_16 = _T_1416;
  assign _T_891_1_17 = _T_1419;
  assign _T_891_1_18 = _T_1422;
  assign _T_891_1_19 = _T_1423;
  assign _T_891_1_20 = _T_1428;
  assign _T_891_1_21 = _T_1431;
  assign _T_891_1_22 = _T_1434;
  assign _T_891_1_23 = _T_1437;
  assign _T_891_1_24 = _T_1440;
  assign _T_891_1_25 = _T_1441;
  assign _T_891_2_0 = _T_1523;
  assign _T_891_2_1 = _T_1524;
  assign _T_891_2_2 = _T_1525;
  assign _T_891_2_3 = _T_1526;
  assign _T_891_2_4 = _T_1527;
  assign _T_891_2_5 = _T_1530;
  assign _T_891_2_6 = _T_1533;
  assign _T_891_2_7 = _T_1536;
  assign _T_891_2_8 = _T_1539;
  assign _T_891_2_9 = _T_1542;
  assign _T_891_2_10 = _T_1543;
  assign _T_891_2_11 = _T_1548;
  assign _T_891_2_12 = _T_1551;
  assign _T_891_2_13 = _T_1554;
  assign _T_891_2_14 = _T_1557;
  assign _T_891_2_15 = _T_1560;
  assign _T_891_2_16 = _T_1563;
  assign _T_891_2_17 = _T_1566;
  assign _T_891_2_18 = _T_1569;
  assign _T_891_2_19 = _T_1570;
  assign _T_891_2_20 = _T_1575;
  assign _T_891_2_21 = _T_1578;
  assign _T_891_2_22 = _T_1581;
  assign _T_891_2_23 = _T_1584;
  assign _T_891_2_24 = _T_1587;
  assign _T_891_2_25 = _T_1588;
  assign ack_back_online = cpu_repair_io_ack_cpus_ok;
  assign cpu_reset_hold_0_io_rst = reset_logic;
  assign cpu_reset_hold_0_io_i = _T_1709;
  assign cpu_reset_hold_1_io_rst = reset_logic;
  assign cpu_reset_hold_1_io_i = _T_1710;
  assign cpu_reset_hold_2_io_rst = reset_logic;
  assign cpu_reset_hold_2_io_i = _T_1711;
  assign reset_all_cpus = cpu_repair_io_reset_cpus;
  assign reset_all_cpus_out = reset_all_cpus_out_hold_io_o;
  assign reset_all_cpus_out_hold_clock = clock;
  assign reset_all_cpus_out_hold_io_rst = reset_logic;
  assign reset_all_cpus_out_hold_io_i = reset_all_cpus;
  assign cpu_repair_io_fault = _T_1972;
  assign cpu_repair_io_cpus_ok = cpu_back_online_reg;
  assign cpu_repair_io_reset_pending = _T_1974;
  assign cpu_repair_io_cpu_in_interrupt = io_cpu_in_interrupt;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_429_aw_ready = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_429_aw_valid = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_429_aw_bits_id = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_429_aw_bits_addr = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_429_aw_bits_len = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_429_aw_bits_size = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_429_aw_bits_burst = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_429_aw_bits_lock = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_429_aw_bits_cache = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_429_aw_bits_prot = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_429_aw_bits_qos = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_429_w_ready = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_429_w_valid = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_429_w_bits_data = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_429_w_bits_strb = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_429_w_bits_last = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_429_b_ready = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  _T_429_b_valid = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  _T_429_b_bits_id = _RAND_18[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  _T_429_b_bits_resp = _RAND_19[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  _T_429_ar_ready = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  _T_429_ar_valid = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  _T_429_ar_bits_id = _RAND_22[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  _T_429_ar_bits_addr = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  _T_429_ar_bits_len = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  _T_429_ar_bits_size = _RAND_25[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  _T_429_ar_bits_burst = _RAND_26[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  _T_429_ar_bits_lock = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  _T_429_ar_bits_cache = _RAND_28[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  _T_429_ar_bits_prot = _RAND_29[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  _T_429_ar_bits_qos = _RAND_30[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  _T_429_r_ready = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  _T_429_r_valid = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  _T_429_r_bits_id = _RAND_33[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  _T_429_r_bits_data = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  _T_429_r_bits_resp = _RAND_35[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  _T_429_r_bits_last = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  _T_487_aw_ready = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  _T_487_aw_valid = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  _T_487_aw_bits_id = _RAND_39[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  _T_487_aw_bits_addr = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  _T_487_aw_bits_len = _RAND_41[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  _T_487_aw_bits_size = _RAND_42[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  _T_487_aw_bits_burst = _RAND_43[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  _T_487_aw_bits_lock = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  _T_487_aw_bits_cache = _RAND_45[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  _T_487_aw_bits_prot = _RAND_46[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  _T_487_aw_bits_qos = _RAND_47[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  _T_487_w_ready = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  _T_487_w_valid = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  _T_487_w_bits_data = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  _T_487_w_bits_strb = _RAND_51[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  _T_487_w_bits_last = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  _T_487_b_ready = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  _T_487_b_valid = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  _T_487_b_bits_id = _RAND_55[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  _T_487_b_bits_resp = _RAND_56[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  _T_487_ar_ready = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  _T_487_ar_valid = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  _T_487_ar_bits_id = _RAND_59[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  _T_487_ar_bits_addr = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  _T_487_ar_bits_len = _RAND_61[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  _T_487_ar_bits_size = _RAND_62[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  _T_487_ar_bits_burst = _RAND_63[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  _T_487_ar_bits_lock = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  _T_487_ar_bits_cache = _RAND_65[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  _T_487_ar_bits_prot = _RAND_66[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  _T_487_ar_bits_qos = _RAND_67[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  _T_487_r_ready = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  _T_487_r_valid = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  _T_487_r_bits_id = _RAND_70[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  _T_487_r_bits_data = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  _T_487_r_bits_resp = _RAND_72[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  _T_487_r_bits_last = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  _T_545_aw_ready = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  _T_545_aw_valid = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  _T_545_aw_bits_id = _RAND_76[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  _T_545_aw_bits_addr = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  _T_545_aw_bits_len = _RAND_78[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  _T_545_aw_bits_size = _RAND_79[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  _T_545_aw_bits_burst = _RAND_80[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  _T_545_aw_bits_lock = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  _T_545_aw_bits_cache = _RAND_82[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  _T_545_aw_bits_prot = _RAND_83[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  _T_545_aw_bits_qos = _RAND_84[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  _T_545_w_ready = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  _T_545_w_valid = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{$random}};
  _T_545_w_bits_data = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{$random}};
  _T_545_w_bits_strb = _RAND_88[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{$random}};
  _T_545_w_bits_last = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{$random}};
  _T_545_b_ready = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{$random}};
  _T_545_b_valid = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{$random}};
  _T_545_b_bits_id = _RAND_92[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{$random}};
  _T_545_b_bits_resp = _RAND_93[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{$random}};
  _T_545_ar_ready = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{$random}};
  _T_545_ar_valid = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{$random}};
  _T_545_ar_bits_id = _RAND_96[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{$random}};
  _T_545_ar_bits_addr = _RAND_97[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{$random}};
  _T_545_ar_bits_len = _RAND_98[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{$random}};
  _T_545_ar_bits_size = _RAND_99[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{$random}};
  _T_545_ar_bits_burst = _RAND_100[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{$random}};
  _T_545_ar_bits_lock = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{$random}};
  _T_545_ar_bits_cache = _RAND_102[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{$random}};
  _T_545_ar_bits_prot = _RAND_103[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{$random}};
  _T_545_ar_bits_qos = _RAND_104[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{$random}};
  _T_545_r_ready = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{$random}};
  _T_545_r_valid = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{$random}};
  _T_545_r_bits_id = _RAND_107[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{$random}};
  _T_545_r_bits_data = _RAND_108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{$random}};
  _T_545_r_bits_resp = _RAND_109[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{$random}};
  _T_545_r_bits_last = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{$random}};
  _T_603_aw_ready = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{$random}};
  _T_603_aw_valid = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{$random}};
  _T_603_aw_bits_id = _RAND_113[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{$random}};
  _T_603_aw_bits_addr = _RAND_114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{$random}};
  _T_603_aw_bits_len = _RAND_115[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{$random}};
  _T_603_aw_bits_size = _RAND_116[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{$random}};
  _T_603_aw_bits_burst = _RAND_117[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{$random}};
  _T_603_aw_bits_lock = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{$random}};
  _T_603_aw_bits_cache = _RAND_119[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{$random}};
  _T_603_aw_bits_prot = _RAND_120[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{$random}};
  _T_603_aw_bits_qos = _RAND_121[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{$random}};
  _T_603_w_ready = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{$random}};
  _T_603_w_valid = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{$random}};
  _T_603_w_bits_data = _RAND_124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{$random}};
  _T_603_w_bits_strb = _RAND_125[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{$random}};
  _T_603_w_bits_last = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{$random}};
  _T_603_b_ready = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{$random}};
  _T_603_b_valid = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{$random}};
  _T_603_b_bits_id = _RAND_129[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{$random}};
  _T_603_b_bits_resp = _RAND_130[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{$random}};
  _T_603_ar_ready = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{$random}};
  _T_603_ar_valid = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{$random}};
  _T_603_ar_bits_id = _RAND_133[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{$random}};
  _T_603_ar_bits_addr = _RAND_134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{$random}};
  _T_603_ar_bits_len = _RAND_135[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{$random}};
  _T_603_ar_bits_size = _RAND_136[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{$random}};
  _T_603_ar_bits_burst = _RAND_137[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{$random}};
  _T_603_ar_bits_lock = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{$random}};
  _T_603_ar_bits_cache = _RAND_139[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{$random}};
  _T_603_ar_bits_prot = _RAND_140[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{$random}};
  _T_603_ar_bits_qos = _RAND_141[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{$random}};
  _T_603_r_ready = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{$random}};
  _T_603_r_valid = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{$random}};
  _T_603_r_bits_id = _RAND_144[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{$random}};
  _T_603_r_bits_data = _RAND_145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{$random}};
  _T_603_r_bits_resp = _RAND_146[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{$random}};
  _T_603_r_bits_last = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{$random}};
  _T_661_aw_ready = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{$random}};
  _T_661_aw_valid = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{$random}};
  _T_661_aw_bits_id = _RAND_150[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{$random}};
  _T_661_aw_bits_addr = _RAND_151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{$random}};
  _T_661_aw_bits_len = _RAND_152[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{$random}};
  _T_661_aw_bits_size = _RAND_153[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{$random}};
  _T_661_aw_bits_burst = _RAND_154[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{$random}};
  _T_661_aw_bits_lock = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{$random}};
  _T_661_aw_bits_cache = _RAND_156[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{$random}};
  _T_661_aw_bits_prot = _RAND_157[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{$random}};
  _T_661_aw_bits_qos = _RAND_158[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{$random}};
  _T_661_w_ready = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{$random}};
  _T_661_w_valid = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{$random}};
  _T_661_w_bits_data = _RAND_161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{$random}};
  _T_661_w_bits_strb = _RAND_162[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{$random}};
  _T_661_w_bits_last = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{$random}};
  _T_661_b_ready = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{$random}};
  _T_661_b_valid = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{$random}};
  _T_661_b_bits_id = _RAND_166[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{$random}};
  _T_661_b_bits_resp = _RAND_167[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{$random}};
  _T_661_ar_ready = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{$random}};
  _T_661_ar_valid = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{$random}};
  _T_661_ar_bits_id = _RAND_170[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{$random}};
  _T_661_ar_bits_addr = _RAND_171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{$random}};
  _T_661_ar_bits_len = _RAND_172[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{$random}};
  _T_661_ar_bits_size = _RAND_173[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{$random}};
  _T_661_ar_bits_burst = _RAND_174[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{$random}};
  _T_661_ar_bits_lock = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{$random}};
  _T_661_ar_bits_cache = _RAND_176[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{$random}};
  _T_661_ar_bits_prot = _RAND_177[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{$random}};
  _T_661_ar_bits_qos = _RAND_178[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{$random}};
  _T_661_r_ready = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{$random}};
  _T_661_r_valid = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{$random}};
  _T_661_r_bits_id = _RAND_181[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{$random}};
  _T_661_r_bits_data = _RAND_182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{$random}};
  _T_661_r_bits_resp = _RAND_183[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{$random}};
  _T_661_r_bits_last = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{$random}};
  _T_719_aw_ready = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{$random}};
  _T_719_aw_valid = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{$random}};
  _T_719_aw_bits_id = _RAND_187[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{$random}};
  _T_719_aw_bits_addr = _RAND_188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{$random}};
  _T_719_aw_bits_len = _RAND_189[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{$random}};
  _T_719_aw_bits_size = _RAND_190[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{$random}};
  _T_719_aw_bits_burst = _RAND_191[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{$random}};
  _T_719_aw_bits_lock = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{$random}};
  _T_719_aw_bits_cache = _RAND_193[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{$random}};
  _T_719_aw_bits_prot = _RAND_194[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{$random}};
  _T_719_aw_bits_qos = _RAND_195[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{$random}};
  _T_719_w_ready = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{$random}};
  _T_719_w_valid = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{$random}};
  _T_719_w_bits_data = _RAND_198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{$random}};
  _T_719_w_bits_strb = _RAND_199[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{$random}};
  _T_719_w_bits_last = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{$random}};
  _T_719_b_ready = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{$random}};
  _T_719_b_valid = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{$random}};
  _T_719_b_bits_id = _RAND_203[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{$random}};
  _T_719_b_bits_resp = _RAND_204[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{$random}};
  _T_719_ar_ready = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{$random}};
  _T_719_ar_valid = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{$random}};
  _T_719_ar_bits_id = _RAND_207[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{$random}};
  _T_719_ar_bits_addr = _RAND_208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{$random}};
  _T_719_ar_bits_len = _RAND_209[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{$random}};
  _T_719_ar_bits_size = _RAND_210[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{$random}};
  _T_719_ar_bits_burst = _RAND_211[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{$random}};
  _T_719_ar_bits_lock = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{$random}};
  _T_719_ar_bits_cache = _RAND_213[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{$random}};
  _T_719_ar_bits_prot = _RAND_214[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{$random}};
  _T_719_ar_bits_qos = _RAND_215[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{$random}};
  _T_719_r_ready = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{$random}};
  _T_719_r_valid = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{$random}};
  _T_719_r_bits_id = _RAND_218[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{$random}};
  _T_719_r_bits_data = _RAND_219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{$random}};
  _T_719_r_bits_resp = _RAND_220[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{$random}};
  _T_719_r_bits_last = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{$random}};
  cpu_reset_im = _RAND_222[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{$random}};
  invalid_reg = _RAND_223[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{$random}};
  faulty_cpu = _RAND_224[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{$random}};
  reset_logic_reg = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{$random}};
  cpu_back_online_reg = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_1713) begin
      _T_429_aw_ready <= _T_487_aw_ready;
    end
    _T_429_aw_valid <= io_cpu0_axi4_aw_valid;
    _T_429_aw_bits_id <= io_cpu0_axi4_aw_bits_id;
    _T_429_aw_bits_addr <= io_cpu0_axi4_aw_bits_addr;
    _T_429_aw_bits_len <= io_cpu0_axi4_aw_bits_len;
    _T_429_aw_bits_size <= io_cpu0_axi4_aw_bits_size;
    _T_429_aw_bits_burst <= io_cpu0_axi4_aw_bits_burst;
    _T_429_aw_bits_lock <= io_cpu0_axi4_aw_bits_lock;
    _T_429_aw_bits_cache <= io_cpu0_axi4_aw_bits_cache;
    _T_429_aw_bits_prot <= io_cpu0_axi4_aw_bits_prot;
    _T_429_aw_bits_qos <= io_cpu0_axi4_aw_bits_qos;
    if (_T_1713) begin
      _T_429_w_ready <= _T_487_w_ready;
    end
    _T_429_w_valid <= io_cpu0_axi4_w_valid;
    _T_429_w_bits_data <= io_cpu0_axi4_w_bits_data;
    _T_429_w_bits_strb <= io_cpu0_axi4_w_bits_strb;
    _T_429_w_bits_last <= io_cpu0_axi4_w_bits_last;
    _T_429_b_ready <= io_cpu0_axi4_b_ready;
    if (_T_1713) begin
      _T_429_b_valid <= _T_487_b_valid;
    end
    if (_T_1713) begin
      _T_429_b_bits_id <= _T_487_b_bits_id;
    end
    if (_T_1713) begin
      _T_429_b_bits_resp <= _T_487_b_bits_resp;
    end
    if (_T_1713) begin
      _T_429_ar_ready <= _T_487_ar_ready;
    end
    _T_429_ar_valid <= io_cpu0_axi4_ar_valid;
    _T_429_ar_bits_id <= io_cpu0_axi4_ar_bits_id;
    _T_429_ar_bits_addr <= io_cpu0_axi4_ar_bits_addr;
    _T_429_ar_bits_len <= io_cpu0_axi4_ar_bits_len;
    _T_429_ar_bits_size <= io_cpu0_axi4_ar_bits_size;
    _T_429_ar_bits_burst <= io_cpu0_axi4_ar_bits_burst;
    _T_429_ar_bits_lock <= io_cpu0_axi4_ar_bits_lock;
    _T_429_ar_bits_cache <= io_cpu0_axi4_ar_bits_cache;
    _T_429_ar_bits_prot <= io_cpu0_axi4_ar_bits_prot;
    _T_429_ar_bits_qos <= io_cpu0_axi4_ar_bits_qos;
    _T_429_r_ready <= io_cpu0_axi4_r_ready;
    if (_T_1713) begin
      _T_429_r_valid <= _T_487_r_valid;
    end
    if (_T_1713) begin
      _T_429_r_bits_id <= _T_487_r_bits_id;
    end
    if (_T_1713) begin
      _T_429_r_bits_data <= _T_487_r_bits_data;
    end
    if (_T_1713) begin
      _T_429_r_bits_resp <= _T_487_r_bits_resp;
    end
    if (_T_1713) begin
      _T_429_r_bits_last <= _T_487_r_bits_last;
    end
    _T_487_aw_ready <= axiBusInternal0_aw_ready;
    if (_T_1713) begin
      _T_487_aw_valid <= _T_429_aw_valid;
    end
    if (_T_1713) begin
      _T_487_aw_bits_id <= _T_429_aw_bits_id;
    end
    if (_T_1713) begin
      _T_487_aw_bits_addr <= _T_429_aw_bits_addr;
    end
    if (_T_1713) begin
      _T_487_aw_bits_len <= _T_429_aw_bits_len;
    end
    if (_T_1713) begin
      _T_487_aw_bits_size <= _T_429_aw_bits_size;
    end
    if (_T_1713) begin
      _T_487_aw_bits_burst <= _T_429_aw_bits_burst;
    end
    if (_T_1713) begin
      _T_487_aw_bits_lock <= _T_429_aw_bits_lock;
    end
    if (_T_1713) begin
      _T_487_aw_bits_cache <= _T_429_aw_bits_cache;
    end
    if (_T_1713) begin
      _T_487_aw_bits_prot <= _T_429_aw_bits_prot;
    end
    if (_T_1713) begin
      _T_487_aw_bits_qos <= _T_429_aw_bits_qos;
    end
    _T_487_w_ready <= axiBusInternal0_w_ready;
    if (_T_1713) begin
      _T_487_w_valid <= _T_429_w_valid;
    end
    if (_T_1713) begin
      _T_487_w_bits_data <= _T_429_w_bits_data;
    end
    if (_T_1713) begin
      _T_487_w_bits_strb <= _T_429_w_bits_strb;
    end
    if (_T_1713) begin
      _T_487_w_bits_last <= _T_429_w_bits_last;
    end
    if (_T_1713) begin
      _T_487_b_ready <= _T_429_b_ready;
    end
    _T_487_b_valid <= axiBusInternal0_b_valid;
    _T_487_b_bits_id <= axiBusInternal0_b_bits_id;
    _T_487_b_bits_resp <= axiBusInternal0_b_bits_resp;
    _T_487_ar_ready <= axiBusInternal0_ar_ready;
    if (_T_1713) begin
      _T_487_ar_valid <= _T_429_ar_valid;
    end
    if (_T_1713) begin
      _T_487_ar_bits_id <= _T_429_ar_bits_id;
    end
    if (_T_1713) begin
      _T_487_ar_bits_addr <= _T_429_ar_bits_addr;
    end
    if (_T_1713) begin
      _T_487_ar_bits_len <= _T_429_ar_bits_len;
    end
    if (_T_1713) begin
      _T_487_ar_bits_size <= _T_429_ar_bits_size;
    end
    if (_T_1713) begin
      _T_487_ar_bits_burst <= _T_429_ar_bits_burst;
    end
    if (_T_1713) begin
      _T_487_ar_bits_lock <= _T_429_ar_bits_lock;
    end
    if (_T_1713) begin
      _T_487_ar_bits_cache <= _T_429_ar_bits_cache;
    end
    if (_T_1713) begin
      _T_487_ar_bits_prot <= _T_429_ar_bits_prot;
    end
    if (_T_1713) begin
      _T_487_ar_bits_qos <= _T_429_ar_bits_qos;
    end
    if (_T_1713) begin
      _T_487_r_ready <= _T_429_r_ready;
    end
    _T_487_r_valid <= axiBusInternal0_r_valid;
    _T_487_r_bits_id <= axiBusInternal0_r_bits_id;
    _T_487_r_bits_data <= axiBusInternal0_r_bits_data;
    _T_487_r_bits_resp <= axiBusInternal0_r_bits_resp;
    _T_487_r_bits_last <= axiBusInternal0_r_bits_last;
    if (_T_1726) begin
      _T_545_aw_ready <= _T_603_aw_ready;
    end
    _T_545_aw_valid <= io_cpu1_axi4_aw_valid;
    _T_545_aw_bits_id <= io_cpu1_axi4_aw_bits_id;
    _T_545_aw_bits_addr <= io_cpu1_axi4_aw_bits_addr;
    _T_545_aw_bits_len <= io_cpu1_axi4_aw_bits_len;
    _T_545_aw_bits_size <= io_cpu1_axi4_aw_bits_size;
    _T_545_aw_bits_burst <= io_cpu1_axi4_aw_bits_burst;
    _T_545_aw_bits_lock <= io_cpu1_axi4_aw_bits_lock;
    _T_545_aw_bits_cache <= io_cpu1_axi4_aw_bits_cache;
    _T_545_aw_bits_prot <= io_cpu1_axi4_aw_bits_prot;
    _T_545_aw_bits_qos <= io_cpu1_axi4_aw_bits_qos;
    if (_T_1726) begin
      _T_545_w_ready <= _T_603_w_ready;
    end
    _T_545_w_valid <= io_cpu1_axi4_w_valid;
    _T_545_w_bits_data <= io_cpu1_axi4_w_bits_data;
    _T_545_w_bits_strb <= io_cpu1_axi4_w_bits_strb;
    _T_545_w_bits_last <= io_cpu1_axi4_w_bits_last;
    _T_545_b_ready <= io_cpu1_axi4_b_ready;
    if (_T_1726) begin
      _T_545_b_valid <= _T_603_b_valid;
    end
    if (_T_1726) begin
      _T_545_b_bits_id <= _T_603_b_bits_id;
    end
    if (_T_1726) begin
      _T_545_b_bits_resp <= _T_603_b_bits_resp;
    end
    if (_T_1726) begin
      _T_545_ar_ready <= _T_603_ar_ready;
    end
    _T_545_ar_valid <= io_cpu1_axi4_ar_valid;
    _T_545_ar_bits_id <= io_cpu1_axi4_ar_bits_id;
    _T_545_ar_bits_addr <= io_cpu1_axi4_ar_bits_addr;
    _T_545_ar_bits_len <= io_cpu1_axi4_ar_bits_len;
    _T_545_ar_bits_size <= io_cpu1_axi4_ar_bits_size;
    _T_545_ar_bits_burst <= io_cpu1_axi4_ar_bits_burst;
    _T_545_ar_bits_lock <= io_cpu1_axi4_ar_bits_lock;
    _T_545_ar_bits_cache <= io_cpu1_axi4_ar_bits_cache;
    _T_545_ar_bits_prot <= io_cpu1_axi4_ar_bits_prot;
    _T_545_ar_bits_qos <= io_cpu1_axi4_ar_bits_qos;
    _T_545_r_ready <= io_cpu1_axi4_r_ready;
    if (_T_1726) begin
      _T_545_r_valid <= _T_603_r_valid;
    end
    if (_T_1726) begin
      _T_545_r_bits_id <= _T_603_r_bits_id;
    end
    if (_T_1726) begin
      _T_545_r_bits_data <= _T_603_r_bits_data;
    end
    if (_T_1726) begin
      _T_545_r_bits_resp <= _T_603_r_bits_resp;
    end
    if (_T_1726) begin
      _T_545_r_bits_last <= _T_603_r_bits_last;
    end
    _T_603_aw_ready <= axiBusInternal1_aw_ready;
    if (_T_1726) begin
      _T_603_aw_valid <= _T_545_aw_valid;
    end
    if (_T_1726) begin
      _T_603_aw_bits_id <= _T_545_aw_bits_id;
    end
    if (_T_1726) begin
      _T_603_aw_bits_addr <= _T_545_aw_bits_addr;
    end
    if (_T_1726) begin
      _T_603_aw_bits_len <= _T_545_aw_bits_len;
    end
    if (_T_1726) begin
      _T_603_aw_bits_size <= _T_545_aw_bits_size;
    end
    if (_T_1726) begin
      _T_603_aw_bits_burst <= _T_545_aw_bits_burst;
    end
    if (_T_1726) begin
      _T_603_aw_bits_lock <= _T_545_aw_bits_lock;
    end
    if (_T_1726) begin
      _T_603_aw_bits_cache <= _T_545_aw_bits_cache;
    end
    if (_T_1726) begin
      _T_603_aw_bits_prot <= _T_545_aw_bits_prot;
    end
    if (_T_1726) begin
      _T_603_aw_bits_qos <= _T_545_aw_bits_qos;
    end
    _T_603_w_ready <= axiBusInternal1_w_ready;
    if (_T_1726) begin
      _T_603_w_valid <= _T_545_w_valid;
    end
    if (_T_1726) begin
      _T_603_w_bits_data <= _T_545_w_bits_data;
    end
    if (_T_1726) begin
      _T_603_w_bits_strb <= _T_545_w_bits_strb;
    end
    if (_T_1726) begin
      _T_603_w_bits_last <= _T_545_w_bits_last;
    end
    if (_T_1726) begin
      _T_603_b_ready <= _T_545_b_ready;
    end
    _T_603_b_valid <= axiBusInternal1_b_valid;
    _T_603_b_bits_id <= axiBusInternal1_b_bits_id;
    _T_603_b_bits_resp <= axiBusInternal1_b_bits_resp;
    _T_603_ar_ready <= axiBusInternal1_ar_ready;
    if (_T_1726) begin
      _T_603_ar_valid <= _T_545_ar_valid;
    end
    if (_T_1726) begin
      _T_603_ar_bits_id <= _T_545_ar_bits_id;
    end
    if (_T_1726) begin
      _T_603_ar_bits_addr <= _T_545_ar_bits_addr;
    end
    if (_T_1726) begin
      _T_603_ar_bits_len <= _T_545_ar_bits_len;
    end
    if (_T_1726) begin
      _T_603_ar_bits_size <= _T_545_ar_bits_size;
    end
    if (_T_1726) begin
      _T_603_ar_bits_burst <= _T_545_ar_bits_burst;
    end
    if (_T_1726) begin
      _T_603_ar_bits_lock <= _T_545_ar_bits_lock;
    end
    if (_T_1726) begin
      _T_603_ar_bits_cache <= _T_545_ar_bits_cache;
    end
    if (_T_1726) begin
      _T_603_ar_bits_prot <= _T_545_ar_bits_prot;
    end
    if (_T_1726) begin
      _T_603_ar_bits_qos <= _T_545_ar_bits_qos;
    end
    if (_T_1726) begin
      _T_603_r_ready <= _T_545_r_ready;
    end
    _T_603_r_valid <= axiBusInternal1_r_valid;
    _T_603_r_bits_id <= axiBusInternal1_r_bits_id;
    _T_603_r_bits_data <= axiBusInternal1_r_bits_data;
    _T_603_r_bits_resp <= axiBusInternal1_r_bits_resp;
    _T_603_r_bits_last <= axiBusInternal1_r_bits_last;
    if (_T_1739) begin
      _T_661_aw_ready <= _T_719_aw_ready;
    end
    _T_661_aw_valid <= io_cpu2_axi4_aw_valid;
    _T_661_aw_bits_id <= io_cpu2_axi4_aw_bits_id;
    _T_661_aw_bits_addr <= io_cpu2_axi4_aw_bits_addr;
    _T_661_aw_bits_len <= io_cpu2_axi4_aw_bits_len;
    _T_661_aw_bits_size <= io_cpu2_axi4_aw_bits_size;
    _T_661_aw_bits_burst <= io_cpu2_axi4_aw_bits_burst;
    _T_661_aw_bits_lock <= io_cpu2_axi4_aw_bits_lock;
    _T_661_aw_bits_cache <= io_cpu2_axi4_aw_bits_cache;
    _T_661_aw_bits_prot <= io_cpu2_axi4_aw_bits_prot;
    _T_661_aw_bits_qos <= io_cpu2_axi4_aw_bits_qos;
    if (_T_1739) begin
      _T_661_w_ready <= _T_719_w_ready;
    end
    _T_661_w_valid <= io_cpu2_axi4_w_valid;
    _T_661_w_bits_data <= io_cpu2_axi4_w_bits_data;
    _T_661_w_bits_strb <= io_cpu2_axi4_w_bits_strb;
    _T_661_w_bits_last <= io_cpu2_axi4_w_bits_last;
    _T_661_b_ready <= io_cpu2_axi4_b_ready;
    if (_T_1739) begin
      _T_661_b_valid <= _T_719_b_valid;
    end
    if (_T_1739) begin
      _T_661_b_bits_id <= _T_719_b_bits_id;
    end
    if (_T_1739) begin
      _T_661_b_bits_resp <= _T_719_b_bits_resp;
    end
    if (_T_1739) begin
      _T_661_ar_ready <= _T_719_ar_ready;
    end
    _T_661_ar_valid <= io_cpu2_axi4_ar_valid;
    _T_661_ar_bits_id <= io_cpu2_axi4_ar_bits_id;
    _T_661_ar_bits_addr <= io_cpu2_axi4_ar_bits_addr;
    _T_661_ar_bits_len <= io_cpu2_axi4_ar_bits_len;
    _T_661_ar_bits_size <= io_cpu2_axi4_ar_bits_size;
    _T_661_ar_bits_burst <= io_cpu2_axi4_ar_bits_burst;
    _T_661_ar_bits_lock <= io_cpu2_axi4_ar_bits_lock;
    _T_661_ar_bits_cache <= io_cpu2_axi4_ar_bits_cache;
    _T_661_ar_bits_prot <= io_cpu2_axi4_ar_bits_prot;
    _T_661_ar_bits_qos <= io_cpu2_axi4_ar_bits_qos;
    _T_661_r_ready <= io_cpu2_axi4_r_ready;
    if (_T_1739) begin
      _T_661_r_valid <= _T_719_r_valid;
    end
    if (_T_1739) begin
      _T_661_r_bits_id <= _T_719_r_bits_id;
    end
    if (_T_1739) begin
      _T_661_r_bits_data <= _T_719_r_bits_data;
    end
    if (_T_1739) begin
      _T_661_r_bits_resp <= _T_719_r_bits_resp;
    end
    if (_T_1739) begin
      _T_661_r_bits_last <= _T_719_r_bits_last;
    end
    _T_719_aw_ready <= axiBusInternal2_aw_ready;
    if (_T_1739) begin
      _T_719_aw_valid <= _T_661_aw_valid;
    end
    if (_T_1739) begin
      _T_719_aw_bits_id <= _T_661_aw_bits_id;
    end
    if (_T_1739) begin
      _T_719_aw_bits_addr <= _T_661_aw_bits_addr;
    end
    if (_T_1739) begin
      _T_719_aw_bits_len <= _T_661_aw_bits_len;
    end
    if (_T_1739) begin
      _T_719_aw_bits_size <= _T_661_aw_bits_size;
    end
    if (_T_1739) begin
      _T_719_aw_bits_burst <= _T_661_aw_bits_burst;
    end
    if (_T_1739) begin
      _T_719_aw_bits_lock <= _T_661_aw_bits_lock;
    end
    if (_T_1739) begin
      _T_719_aw_bits_cache <= _T_661_aw_bits_cache;
    end
    if (_T_1739) begin
      _T_719_aw_bits_prot <= _T_661_aw_bits_prot;
    end
    if (_T_1739) begin
      _T_719_aw_bits_qos <= _T_661_aw_bits_qos;
    end
    _T_719_w_ready <= axiBusInternal2_w_ready;
    if (_T_1739) begin
      _T_719_w_valid <= _T_661_w_valid;
    end
    if (_T_1739) begin
      _T_719_w_bits_data <= _T_661_w_bits_data;
    end
    if (_T_1739) begin
      _T_719_w_bits_strb <= _T_661_w_bits_strb;
    end
    if (_T_1739) begin
      _T_719_w_bits_last <= _T_661_w_bits_last;
    end
    if (_T_1739) begin
      _T_719_b_ready <= _T_661_b_ready;
    end
    _T_719_b_valid <= axiBusInternal2_b_valid;
    _T_719_b_bits_id <= axiBusInternal2_b_bits_id;
    _T_719_b_bits_resp <= axiBusInternal2_b_bits_resp;
    _T_719_ar_ready <= axiBusInternal2_ar_ready;
    if (_T_1739) begin
      _T_719_ar_valid <= _T_661_ar_valid;
    end
    if (_T_1739) begin
      _T_719_ar_bits_id <= _T_661_ar_bits_id;
    end
    if (_T_1739) begin
      _T_719_ar_bits_addr <= _T_661_ar_bits_addr;
    end
    if (_T_1739) begin
      _T_719_ar_bits_len <= _T_661_ar_bits_len;
    end
    if (_T_1739) begin
      _T_719_ar_bits_size <= _T_661_ar_bits_size;
    end
    if (_T_1739) begin
      _T_719_ar_bits_burst <= _T_661_ar_bits_burst;
    end
    if (_T_1739) begin
      _T_719_ar_bits_lock <= _T_661_ar_bits_lock;
    end
    if (_T_1739) begin
      _T_719_ar_bits_cache <= _T_661_ar_bits_cache;
    end
    if (_T_1739) begin
      _T_719_ar_bits_prot <= _T_661_ar_bits_prot;
    end
    if (_T_1739) begin
      _T_719_ar_bits_qos <= _T_661_ar_bits_qos;
    end
    if (_T_1739) begin
      _T_719_r_ready <= _T_661_r_ready;
    end
    _T_719_r_valid <= axiBusInternal2_r_valid;
    _T_719_r_bits_id <= axiBusInternal2_r_bits_id;
    _T_719_r_bits_data <= axiBusInternal2_r_bits_data;
    _T_719_r_bits_resp <= axiBusInternal2_r_bits_resp;
    _T_719_r_bits_last <= axiBusInternal2_r_bits_last;
    if (_T_1704) begin
      cpu_reset_im <= _T_1705;
    end else begin
      cpu_reset_im <= 3'h0;
    end
    if (reset) begin
      invalid_reg <= 3'h0;
    end else begin
      invalid_reg <= _GEN_12[2:0];
    end
    if (reset) begin
      faulty_cpu <= 3'h0;
    end else begin
      if (_T_1704) begin
        faulty_cpu <= _T_1705;
      end else begin
        faulty_cpu <= 3'h0;
      end
    end
    if (reset) begin
      reset_logic_reg <= 1'h0;
    end else begin
      if (reset_logic_reg) begin
        if (_T_1693) begin
          reset_logic_reg <= 1'h0;
        end else begin
          if (reset_logic) begin
            reset_logic_reg <= 1'h1;
          end
        end
      end else begin
        if (reset_logic) begin
          reset_logic_reg <= 1'h1;
        end
      end
    end
    if (reset) begin
      cpu_back_online_reg <= 1'h0;
    end else begin
      if (ack_back_online) begin
        cpu_back_online_reg <= 1'h0;
      end else begin
        if (reset_logic_reg) begin
          if (_T_1693) begin
            cpu_back_online_reg <= 1'h1;
          end
        end
      end
    end
  end
endmodule


`timescale 1 ns / 1 ps

	module fault_detector_v1_0 #
	(

		// Parameters of Axi Slave Bus Interface CPU0_AXI
		parameter integer C_CPU0_AXI_ID_WIDTH	= 4,
		parameter integer C_CPU0_AXI_DATA_WIDTH	= 32,
		parameter integer C_CPU0_AXI_ADDR_WIDTH	= 32,
		parameter integer C_CPU0_AXI_AWUSER_WIDTH	= 0,
		parameter integer C_CPU0_AXI_ARUSER_WIDTH	= 0,
		parameter integer C_CPU0_AXI_WUSER_WIDTH	= 0,
		parameter integer C_CPU0_AXI_RUSER_WIDTH	= 0,
		parameter integer C_CPU0_AXI_BUSER_WIDTH	= 0,

		// Parameters of Axi Slave Bus Interface CPU1_AXI
		parameter integer C_CPU1_AXI_ID_WIDTH	= 4,
		parameter integer C_CPU1_AXI_DATA_WIDTH	= 32,
		parameter integer C_CPU1_AXI_ADDR_WIDTH	= 32,
		parameter integer C_CPU1_AXI_AWUSER_WIDTH	= 0,
		parameter integer C_CPU1_AXI_ARUSER_WIDTH	= 0,
		parameter integer C_CPU1_AXI_WUSER_WIDTH	= 0,
		parameter integer C_CPU1_AXI_RUSER_WIDTH	= 0,
		parameter integer C_CPU1_AXI_BUSER_WIDTH	= 0,

		// Parameters of Axi Slave Bus Interface CPU2_AXI
		parameter integer C_CPU2_AXI_ID_WIDTH	= 4,
		parameter integer C_CPU2_AXI_DATA_WIDTH	= 32,
		parameter integer C_CPU2_AXI_ADDR_WIDTH	= 32,
		parameter integer C_CPU2_AXI_AWUSER_WIDTH	= 0,
		parameter integer C_CPU2_AXI_ARUSER_WIDTH	= 0,
		parameter integer C_CPU2_AXI_WUSER_WIDTH	= 0,
		parameter integer C_CPU2_AXI_RUSER_WIDTH	= 0,
		parameter integer C_CPU2_AXI_BUSER_WIDTH	= 0,

		// Parameters of Axi Master Bus Interface OUT_AXI
		parameter  C_OUT_AXI_TARGET_SLAVE_BASE_ADDR	= 32'h40000000,
		parameter integer C_OUT_AXI_BURST_LEN	= 16,
		parameter integer C_OUT_AXI_ID_WIDTH	= 4,
		parameter integer C_OUT_AXI_ADDR_WIDTH	= 32,
		parameter integer C_OUT_AXI_DATA_WIDTH	= 32,
		parameter integer C_OUT_AXI_AWUSER_WIDTH	= 0,
		parameter integer C_OUT_AXI_ARUSER_WIDTH	= 0,
		parameter integer C_OUT_AXI_WUSER_WIDTH	= 0,
		parameter integer C_OUT_AXI_RUSER_WIDTH	= 0,
		parameter integer C_OUT_AXI_BUSER_WIDTH	= 0
	)
	(

		// Ports of Axi Slave Bus Interface CPU0_AXI
		input wire  cpu0_axi_aclk,
		input wire  cpu0_axi_aresetn,
		input wire [C_CPU0_AXI_ID_WIDTH-1 : 0] cpu0_axi_awid,
		input wire [C_CPU0_AXI_ADDR_WIDTH-1 : 0] cpu0_axi_awaddr,
		input wire [7 : 0] cpu0_axi_awlen,
		input wire [2 : 0] cpu0_axi_awsize,
		input wire [1 : 0] cpu0_axi_awburst,
		input wire  cpu0_axi_awlock,
		input wire [3 : 0] cpu0_axi_awcache,
		input wire [2 : 0] cpu0_axi_awprot,
		input wire [3 : 0] cpu0_axi_awqos,
		input wire [3 : 0] cpu0_axi_awregion,
		input wire [C_CPU0_AXI_AWUSER_WIDTH-1 : 0] cpu0_axi_awuser,
		input wire  cpu0_axi_awvalid,
		output wire  cpu0_axi_awready,
		input wire [C_CPU0_AXI_DATA_WIDTH-1 : 0] cpu0_axi_wdata,
		input wire [(C_CPU0_AXI_DATA_WIDTH/8)-1 : 0] cpu0_axi_wstrb,
		input wire  cpu0_axi_wlast,
		input wire [C_CPU0_AXI_WUSER_WIDTH-1 : 0] cpu0_axi_wuser,
		input wire  cpu0_axi_wvalid,
		output wire  cpu0_axi_wready,
		output wire [C_CPU0_AXI_ID_WIDTH-1 : 0] cpu0_axi_bid,
		output wire [1 : 0] cpu0_axi_bresp,
		output wire [C_CPU0_AXI_BUSER_WIDTH-1 : 0] cpu0_axi_buser,
		output wire  cpu0_axi_bvalid,
		input wire  cpu0_axi_bready,
		input wire [C_CPU0_AXI_ID_WIDTH-1 : 0] cpu0_axi_arid,
		input wire [C_CPU0_AXI_ADDR_WIDTH-1 : 0] cpu0_axi_araddr,
		input wire [7 : 0] cpu0_axi_arlen,
		input wire [2 : 0] cpu0_axi_arsize,
		input wire [1 : 0] cpu0_axi_arburst,
		input wire  cpu0_axi_arlock,
		input wire [3 : 0] cpu0_axi_arcache,
		input wire [2 : 0] cpu0_axi_arprot,
		input wire [3 : 0] cpu0_axi_arqos,
		input wire [3 : 0] cpu0_axi_arregion,
		input wire [C_CPU0_AXI_ARUSER_WIDTH-1 : 0] cpu0_axi_aruser,
		input wire  cpu0_axi_arvalid,
		output wire  cpu0_axi_arready,
		output wire [C_CPU0_AXI_ID_WIDTH-1 : 0] cpu0_axi_rid,
		output wire [C_CPU0_AXI_DATA_WIDTH-1 : 0] cpu0_axi_rdata,
		output wire [1 : 0] cpu0_axi_rresp,
		output wire  cpu0_axi_rlast,
		output wire [C_CPU0_AXI_RUSER_WIDTH-1 : 0] cpu0_axi_ruser,
		output wire  cpu0_axi_rvalid,
		input wire  cpu0_axi_rready,

		// Ports of Axi Slave Bus Interface CPU1_AXI
		input wire  cpu1_axi_aclk,
		input wire  cpu1_axi_aresetn,
		input wire [C_CPU1_AXI_ID_WIDTH-1 : 0] cpu1_axi_awid,
		input wire [C_CPU1_AXI_ADDR_WIDTH-1 : 0] cpu1_axi_awaddr,
		input wire [7 : 0] cpu1_axi_awlen,
		input wire [2 : 0] cpu1_axi_awsize,
		input wire [1 : 0] cpu1_axi_awburst,
		input wire  cpu1_axi_awlock,
		input wire [3 : 0] cpu1_axi_awcache,
		input wire [2 : 0] cpu1_axi_awprot,
		input wire [3 : 0] cpu1_axi_awqos,
		input wire [3 : 0] cpu1_axi_awregion,
		input wire [C_CPU1_AXI_AWUSER_WIDTH-1 : 0] cpu1_axi_awuser,
		input wire  cpu1_axi_awvalid,
		output wire  cpu1_axi_awready,
		input wire [C_CPU1_AXI_DATA_WIDTH-1 : 0] cpu1_axi_wdata,
		input wire [(C_CPU1_AXI_DATA_WIDTH/8)-1 : 0] cpu1_axi_wstrb,
		input wire  cpu1_axi_wlast,
		input wire [C_CPU1_AXI_WUSER_WIDTH-1 : 0] cpu1_axi_wuser,
		input wire  cpu1_axi_wvalid,
		output wire  cpu1_axi_wready,
		output wire [C_CPU1_AXI_ID_WIDTH-1 : 0] cpu1_axi_bid,
		output wire [1 : 0] cpu1_axi_bresp,
		output wire [C_CPU1_AXI_BUSER_WIDTH-1 : 0] cpu1_axi_buser,
		output wire  cpu1_axi_bvalid,
		input wire  cpu1_axi_bready,
		input wire [C_CPU1_AXI_ID_WIDTH-1 : 0] cpu1_axi_arid,
		input wire [C_CPU1_AXI_ADDR_WIDTH-1 : 0] cpu1_axi_araddr,
		input wire [7 : 0] cpu1_axi_arlen,
		input wire [2 : 0] cpu1_axi_arsize,
		input wire [1 : 0] cpu1_axi_arburst,
		input wire  cpu1_axi_arlock,
		input wire [3 : 0] cpu1_axi_arcache,
		input wire [2 : 0] cpu1_axi_arprot,
		input wire [3 : 0] cpu1_axi_arqos,
		input wire [3 : 0] cpu1_axi_arregion,
		input wire [C_CPU1_AXI_ARUSER_WIDTH-1 : 0] cpu1_axi_aruser,
		input wire  cpu1_axi_arvalid,
		output wire  cpu1_axi_arready,
		output wire [C_CPU1_AXI_ID_WIDTH-1 : 0] cpu1_axi_rid,
		output wire [C_CPU1_AXI_DATA_WIDTH-1 : 0] cpu1_axi_rdata,
		output wire [1 : 0] cpu1_axi_rresp,
		output wire  cpu1_axi_rlast,
		output wire [C_CPU1_AXI_RUSER_WIDTH-1 : 0] cpu1_axi_ruser,
		output wire  cpu1_axi_rvalid,
		input wire  cpu1_axi_rready,

		// Ports of Axi Slave Bus Interface CPU2_AXI
		input wire  cpu2_axi_aclk,
		input wire  cpu2_axi_aresetn,
		input wire [C_CPU2_AXI_ID_WIDTH-1 : 0] cpu2_axi_awid,
		input wire [C_CPU2_AXI_ADDR_WIDTH-1 : 0] cpu2_axi_awaddr,
		input wire [7 : 0] cpu2_axi_awlen,
		input wire [2 : 0] cpu2_axi_awsize,
		input wire [1 : 0] cpu2_axi_awburst,
		input wire  cpu2_axi_awlock,
		input wire [3 : 0] cpu2_axi_awcache,
		input wire [2 : 0] cpu2_axi_awprot,
		input wire [3 : 0] cpu2_axi_awqos,
		input wire [3 : 0] cpu2_axi_awregion,
		input wire [C_CPU2_AXI_AWUSER_WIDTH-1 : 0] cpu2_axi_awuser,
		input wire  cpu2_axi_awvalid,
		output wire  cpu2_axi_awready,
		input wire [C_CPU2_AXI_DATA_WIDTH-1 : 0] cpu2_axi_wdata,
		input wire [(C_CPU2_AXI_DATA_WIDTH/8)-1 : 0] cpu2_axi_wstrb,
		input wire  cpu2_axi_wlast,
		input wire [C_CPU2_AXI_WUSER_WIDTH-1 : 0] cpu2_axi_wuser,
		input wire  cpu2_axi_wvalid,
		output wire  cpu2_axi_wready,
		output wire [C_CPU2_AXI_ID_WIDTH-1 : 0] cpu2_axi_bid,
		output wire [1 : 0] cpu2_axi_bresp,
		output wire [C_CPU2_AXI_BUSER_WIDTH-1 : 0] cpu2_axi_buser,
		output wire  cpu2_axi_bvalid,
		input wire  cpu2_axi_bready,
		input wire [C_CPU2_AXI_ID_WIDTH-1 : 0] cpu2_axi_arid,
		input wire [C_CPU2_AXI_ADDR_WIDTH-1 : 0] cpu2_axi_araddr,
		input wire [7 : 0] cpu2_axi_arlen,
		input wire [2 : 0] cpu2_axi_arsize,
		input wire [1 : 0] cpu2_axi_arburst,
		input wire  cpu2_axi_arlock,
		input wire [3 : 0] cpu2_axi_arcache,
		input wire [2 : 0] cpu2_axi_arprot,
		input wire [3 : 0] cpu2_axi_arqos,
		input wire [3 : 0] cpu2_axi_arregion,
		input wire [C_CPU2_AXI_ARUSER_WIDTH-1 : 0] cpu2_axi_aruser,
		input wire  cpu2_axi_arvalid,
		output wire  cpu2_axi_arready,
		output wire [C_CPU2_AXI_ID_WIDTH-1 : 0] cpu2_axi_rid,
		output wire [C_CPU2_AXI_DATA_WIDTH-1 : 0] cpu2_axi_rdata,
		output wire [1 : 0] cpu2_axi_rresp,
		output wire  cpu2_axi_rlast,
		output wire [C_CPU2_AXI_RUSER_WIDTH-1 : 0] cpu2_axi_ruser,
		output wire  cpu2_axi_rvalid,
		input wire  cpu2_axi_rready,

		// Ports of Axi Master Bus Interface OUT_AXI
		input wire  out_axi_aclk,
		input wire  out_axi_aresetn,
		output wire [C_OUT_AXI_ID_WIDTH-1 : 0] out_axi_awid,
		output wire [C_OUT_AXI_ADDR_WIDTH-1 : 0] out_axi_awaddr,
		output wire [7 : 0] out_axi_awlen,
		output wire [2 : 0] out_axi_awsize,
		output wire [1 : 0] out_axi_awburst,
		output wire  out_axi_awlock,
		output wire [3 : 0] out_axi_awcache,
		output wire [2 : 0] out_axi_awprot,
		output wire [3 : 0] out_axi_awqos,
		output wire [C_OUT_AXI_AWUSER_WIDTH-1 : 0] out_axi_awuser,
		output wire  out_axi_awvalid,
		input wire  out_axi_awready,
		output wire [C_OUT_AXI_DATA_WIDTH-1 : 0] out_axi_wdata,
		output wire [C_OUT_AXI_DATA_WIDTH/8-1 : 0] out_axi_wstrb,
		output wire  out_axi_wlast,
		output wire [C_OUT_AXI_WUSER_WIDTH-1 : 0] out_axi_wuser,
		output wire  out_axi_wvalid,
		input wire  out_axi_wready,
		input wire [C_OUT_AXI_ID_WIDTH-1 : 0] out_axi_bid,
		input wire [1 : 0] out_axi_bresp,
		input wire [C_OUT_AXI_BUSER_WIDTH-1 : 0] out_axi_buser,
		input wire  out_axi_bvalid,
		output wire  out_axi_bready,
		output wire [C_OUT_AXI_ID_WIDTH-1 : 0] out_axi_arid,
		output wire [C_OUT_AXI_ADDR_WIDTH-1 : 0] out_axi_araddr,
		output wire [7 : 0] out_axi_arlen,
		output wire [2 : 0] out_axi_arsize,
		output wire [1 : 0] out_axi_arburst,
		output wire  out_axi_arlock,
		output wire [3 : 0] out_axi_arcache,
		output wire [2 : 0] out_axi_arprot,
		output wire [3 : 0] out_axi_arqos,
		output wire [C_OUT_AXI_ARUSER_WIDTH-1 : 0] out_axi_aruser,
		output wire  out_axi_arvalid,
		input wire  out_axi_arready,
		input wire [C_OUT_AXI_ID_WIDTH-1 : 0] out_axi_rid,
		input wire [C_OUT_AXI_DATA_WIDTH-1 : 0] out_axi_rdata,
		input wire [1 : 0] out_axi_rresp,
		input wire  out_axi_rlast,
		input wire [C_OUT_AXI_RUSER_WIDTH-1 : 0] out_axi_ruser,
		input wire  out_axi_rvalid,
		output wire  out_axi_rready,

		output wire [2:0] invalid,
		output wire [2:0] fault_reset_vector,
		output wire [2:0] reset_cpu,
		input wire reset_disable,
		input wire [2:0] reset_routing_logic,
		output wire cpu_back_online,
		input wire ack_back_online,
		output wire stop_all_cpus,
		output wire latch_registers,
		output wire reset_to_recovery,
		input wire cpu_reset_feedback,
		input wire cpu_in_interrupt
	);

    wire reset;
    assign reset = ~(out_axi_aresetn);

	assign out_axi_wuser = 0;
	assign out_axi_aruser = 0;
    assign out_axi_awuser = 0;

	assign cpu0_axi_ruser = 0;
	assign cpu1_axi_ruser = 0;
	assign cpu2_axi_ruser = 0;

	assign cpu0_axi_buser = 0;
	assign cpu1_axi_buser = 0;
	assign cpu2_axi_buser = 0;

    FaultDetector fault_detector_inst (

		.clock(out_axi_aclk),
		.reset(reset),
		.io_invalid(invalid),
		.io_fault_reset_vector(fault_reset_vector),
		.io_reset_cpu(reset_cpu),
		.io_disable_reset(reset_disable),
		.io_reset_routing_logic(reset_routing_logic),
		.io_cpu_back_online(cpu_back_online),
		.io_ack_back_online(ack_back_online),
		.io_stop_all_cpus(stop_all_cpus),
		.io_latch_registers(latch_registers),
		.io_reset_to_recovery(reset_to_recovery),
		.io_cpu_reset_feedback(cpu_reset_feedback),
		.io_cpu_in_interrupt(cpu_in_interrupt),

		.io_cpu0_axi4_aw_ready(cpu0_axi_awready),
		.io_cpu0_axi4_aw_valid(cpu0_axi_awvalid),
		.io_cpu0_axi4_aw_bits_id(cpu0_axi_awid),
		.io_cpu0_axi4_aw_bits_addr(cpu0_axi_awaddr),
		.io_cpu0_axi4_aw_bits_len(cpu0_axi_awlen),
		.io_cpu0_axi4_aw_bits_size(cpu0_axi_awsize),
		.io_cpu0_axi4_aw_bits_burst(cpu0_axi_awburst),
		.io_cpu0_axi4_aw_bits_lock(cpu0_axi_awlock),
		.io_cpu0_axi4_aw_bits_cache(cpu0_axi_awcache),
		.io_cpu0_axi4_aw_bits_prot(cpu0_axi_awprot),
		.io_cpu0_axi4_aw_bits_qos(cpu0_axi_awqos),

		.io_cpu0_axi4_w_ready(cpu0_axi_wready),
		.io_cpu0_axi4_w_valid(cpu0_axi_wvalid),
		.io_cpu0_axi4_w_bits_data(cpu0_axi_wdata),
		.io_cpu0_axi4_w_bits_strb(cpu0_axi_wstrb),
		.io_cpu0_axi4_w_bits_last(cpu0_axi_wlast),

		.io_cpu0_axi4_b_ready(cpu0_axi_bready),
		.io_cpu0_axi4_b_valid(cpu0_axi_bvalid),
		.io_cpu0_axi4_b_bits_id(cpu0_axi_bid),
		.io_cpu0_axi4_b_bits_resp(cpu0_axi_bresp),

		.io_cpu0_axi4_ar_ready(cpu0_axi_arready),
		.io_cpu0_axi4_ar_valid(cpu0_axi_arvalid),
		.io_cpu0_axi4_ar_bits_id(cpu0_axi_arid),
		.io_cpu0_axi4_ar_bits_addr(cpu0_axi_araddr),
		.io_cpu0_axi4_ar_bits_len(cpu0_axi_arlen),
		.io_cpu0_axi4_ar_bits_size(cpu0_axi_arsize),
		.io_cpu0_axi4_ar_bits_burst(cpu0_axi_arburst),
		.io_cpu0_axi4_ar_bits_lock(cpu0_axi_arlock),
		.io_cpu0_axi4_ar_bits_cache(cpu0_axi_arcache),
		.io_cpu0_axi4_ar_bits_prot(cpu0_axi_arprot),
		.io_cpu0_axi4_ar_bits_qos(cpu0_axi_arqos),

		.io_cpu0_axi4_r_ready(cpu0_axi_rready),
		.io_cpu0_axi4_r_valid(cpu0_axi_rvalid),
		.io_cpu0_axi4_r_bits_id(cpu0_axi_rid),
		.io_cpu0_axi4_r_bits_data(cpu0_axi_rdata),
		.io_cpu0_axi4_r_bits_resp(cpu0_axi_rresp),
		.io_cpu0_axi4_r_bits_last(cpu0_axi_rlast),

		// CPU1
		.io_cpu1_axi4_aw_ready(cpu1_axi_awready),
		.io_cpu1_axi4_aw_valid(cpu1_axi_awvalid),
		.io_cpu1_axi4_aw_bits_id(cpu1_axi_awid),
		.io_cpu1_axi4_aw_bits_addr(cpu1_axi_awaddr),
		.io_cpu1_axi4_aw_bits_len(cpu1_axi_awlen),
		.io_cpu1_axi4_aw_bits_size(cpu1_axi_awsize),
		.io_cpu1_axi4_aw_bits_burst(cpu1_axi_awburst),
		.io_cpu1_axi4_aw_bits_lock(cpu1_axi_awlock),
		.io_cpu1_axi4_aw_bits_cache(cpu1_axi_awcache),
		.io_cpu1_axi4_aw_bits_prot(cpu1_axi_awprot),
		.io_cpu1_axi4_aw_bits_qos(cpu1_axi_awqos),

		.io_cpu1_axi4_w_ready(cpu1_axi_wready),
		.io_cpu1_axi4_w_valid(cpu1_axi_wvalid),
		.io_cpu1_axi4_w_bits_data(cpu1_axi_wdata),
		.io_cpu1_axi4_w_bits_strb(cpu1_axi_wstrb),
		.io_cpu1_axi4_w_bits_last(cpu1_axi_wlast),

		.io_cpu1_axi4_b_ready(cpu1_axi_bready),
		.io_cpu1_axi4_b_valid(cpu1_axi_bvalid),
		.io_cpu1_axi4_b_bits_id(cpu1_axi_bid),
		.io_cpu1_axi4_b_bits_resp(cpu1_axi_bresp),

		.io_cpu1_axi4_ar_ready(cpu1_axi_arready),
		.io_cpu1_axi4_ar_valid(cpu1_axi_arvalid),
		.io_cpu1_axi4_ar_bits_id(cpu1_axi_arid),
		.io_cpu1_axi4_ar_bits_addr(cpu1_axi_araddr),
		.io_cpu1_axi4_ar_bits_len(cpu1_axi_arlen),
		.io_cpu1_axi4_ar_bits_size(cpu1_axi_arsize),
		.io_cpu1_axi4_ar_bits_burst(cpu1_axi_arburst),
		.io_cpu1_axi4_ar_bits_lock(cpu1_axi_arlock),
		.io_cpu1_axi4_ar_bits_cache(cpu1_axi_arcache),
		.io_cpu1_axi4_ar_bits_prot(cpu1_axi_arprot),
		.io_cpu1_axi4_ar_bits_qos(cpu1_axi_arqos),

		.io_cpu1_axi4_r_ready(cpu1_axi_rready),
		.io_cpu1_axi4_r_valid(cpu1_axi_rvalid),
		.io_cpu1_axi4_r_bits_id(cpu1_axi_rid),
		.io_cpu1_axi4_r_bits_data(cpu1_axi_rdata),
		.io_cpu1_axi4_r_bits_resp(cpu1_axi_rresp),
		.io_cpu1_axi4_r_bits_last(cpu1_axi_rlast),

		// CPU2
		.io_cpu2_axi4_aw_ready(cpu2_axi_awready),
		.io_cpu2_axi4_aw_valid(cpu2_axi_awvalid),
		.io_cpu2_axi4_aw_bits_id(cpu2_axi_awid),
		.io_cpu2_axi4_aw_bits_addr(cpu2_axi_awaddr),
		.io_cpu2_axi4_aw_bits_len(cpu2_axi_awlen),
		.io_cpu2_axi4_aw_bits_size(cpu2_axi_awsize),
		.io_cpu2_axi4_aw_bits_burst(cpu2_axi_awburst),
		.io_cpu2_axi4_aw_bits_lock(cpu2_axi_awlock),
		.io_cpu2_axi4_aw_bits_cache(cpu2_axi_awcache),
		.io_cpu2_axi4_aw_bits_prot(cpu2_axi_awprot),
		.io_cpu2_axi4_aw_bits_qos(cpu2_axi_awqos),

		.io_cpu2_axi4_w_ready(cpu2_axi_wready),
		.io_cpu2_axi4_w_valid(cpu2_axi_wvalid),
		.io_cpu2_axi4_w_bits_data(cpu2_axi_wdata),
		.io_cpu2_axi4_w_bits_strb(cpu2_axi_wstrb),
		.io_cpu2_axi4_w_bits_last(cpu2_axi_wlast),

		.io_cpu2_axi4_b_ready(cpu2_axi_bready),
		.io_cpu2_axi4_b_valid(cpu2_axi_bvalid),
		.io_cpu2_axi4_b_bits_id(cpu2_axi_bid),
		.io_cpu2_axi4_b_bits_resp(cpu2_axi_bresp),

		.io_cpu2_axi4_ar_ready(cpu2_axi_arready),
		.io_cpu2_axi4_ar_valid(cpu2_axi_arvalid),
		.io_cpu2_axi4_ar_bits_id(cpu2_axi_arid),
		.io_cpu2_axi4_ar_bits_addr(cpu2_axi_araddr),
		.io_cpu2_axi4_ar_bits_len(cpu2_axi_arlen),
		.io_cpu2_axi4_ar_bits_size(cpu2_axi_arsize),
		.io_cpu2_axi4_ar_bits_burst(cpu2_axi_arburst),
		.io_cpu2_axi4_ar_bits_lock(cpu2_axi_arlock),
		.io_cpu2_axi4_ar_bits_cache(cpu2_axi_arcache),
		.io_cpu2_axi4_ar_bits_prot(cpu2_axi_arprot),
		.io_cpu2_axi4_ar_bits_qos(cpu2_axi_arqos),

		.io_cpu2_axi4_r_ready(cpu2_axi_rready),
		.io_cpu2_axi4_r_valid(cpu2_axi_rvalid),
		.io_cpu2_axi4_r_bits_id(cpu2_axi_rid),
		.io_cpu2_axi4_r_bits_data(cpu2_axi_rdata),
		.io_cpu2_axi4_r_bits_resp(cpu2_axi_rresp),
		.io_cpu2_axi4_r_bits_last(cpu2_axi_rlast),

		// OUT
		.io_out_axi4_aw_ready(out_axi_awready),
		.io_out_axi4_aw_valid(out_axi_awvalid),
		.io_out_axi4_aw_bits_id(out_axi_awid),
		.io_out_axi4_aw_bits_addr(out_axi_awaddr),
		.io_out_axi4_aw_bits_len(out_axi_awlen),
		.io_out_axi4_aw_bits_size(out_axi_awsize),
		.io_out_axi4_aw_bits_burst(out_axi_awburst),
		.io_out_axi4_aw_bits_lock(out_axi_awlock),
		.io_out_axi4_aw_bits_cache(out_axi_awcache),
		.io_out_axi4_aw_bits_prot(out_axi_awprot),
		.io_out_axi4_aw_bits_qos(out_axi_awqos),

		.io_out_axi4_w_ready(out_axi_wready),
		.io_out_axi4_w_valid(out_axi_wvalid),
		.io_out_axi4_w_bits_data(out_axi_wdata),
		.io_out_axi4_w_bits_strb(out_axi_wstrb),
		.io_out_axi4_w_bits_last(out_axi_wlast),

		.io_out_axi4_b_ready(out_axi_bready),
		.io_out_axi4_b_valid(out_axi_bvalid),
		.io_out_axi4_b_bits_id(out_axi_bid),
		.io_out_axi4_b_bits_resp(out_axi_bresp),

		.io_out_axi4_ar_ready(out_axi_arready),
		.io_out_axi4_ar_valid(out_axi_arvalid),
		.io_out_axi4_ar_bits_id(out_axi_arid),
		.io_out_axi4_ar_bits_addr(out_axi_araddr),
		.io_out_axi4_ar_bits_len(out_axi_arlen),
		.io_out_axi4_ar_bits_size(out_axi_arsize),
		.io_out_axi4_ar_bits_burst(out_axi_arburst),
		.io_out_axi4_ar_bits_lock(out_axi_arlock),
		.io_out_axi4_ar_bits_cache(out_axi_arcache),
		.io_out_axi4_ar_bits_prot(out_axi_arprot),
		.io_out_axi4_ar_bits_qos(out_axi_arqos),

		.io_out_axi4_r_ready(out_axi_rready),
		.io_out_axi4_r_valid(out_axi_rvalid),
		.io_out_axi4_r_bits_id(out_axi_rid),
		.io_out_axi4_r_bits_data(out_axi_rdata),
		.io_out_axi4_r_bits_resp(out_axi_rresp),
		.io_out_axi4_r_bits_last(out_axi_rlast)
	);


	endmodule
